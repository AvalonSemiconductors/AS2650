module ram_controller (CEN_all,
    GWEN_0,
    GWEN_1,
    GWEN_2,
    GWEN_3,
    GWEN_4,
    GWEN_5,
    GWEN_6,
    GWEN_7,
    WEb_ram,
    ram_enabled,
    rst,
    vdd,
    vss,
    wb_clk_i,
    A_all,
    D_all,
    Q0,
    Q1,
    Q2,
    Q3,
    Q4,
    Q5,
    Q6,
    Q7,
    WEN_all,
    bus_in,
    bus_out,
    requested_addr);
 output CEN_all;
 output GWEN_0;
 output GWEN_1;
 output GWEN_2;
 output GWEN_3;
 output GWEN_4;
 output GWEN_5;
 output GWEN_6;
 output GWEN_7;
 input WEb_ram;
 input ram_enabled;
 input rst;
 input vdd;
 input vss;
 input wb_clk_i;
 output [8:0] A_all;
 output [7:0] D_all;
 input [7:0] Q0;
 input [7:0] Q1;
 input [7:0] Q2;
 input [7:0] Q3;
 input [7:0] Q4;
 input [7:0] Q5;
 input [7:0] Q6;
 input [7:0] Q7;
 output [7:0] WEN_all;
 input [7:0] bus_in;
 output [7:0] bus_out;
 input [15:0] requested_addr;

 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \requested_addr_latch[0] ;
 wire \requested_addr_latch[10] ;
 wire \requested_addr_latch[11] ;
 wire \requested_addr_latch[12] ;
 wire \requested_addr_latch[13] ;
 wire \requested_addr_latch[14] ;
 wire \requested_addr_latch[15] ;
 wire \requested_addr_latch[1] ;
 wire \requested_addr_latch[2] ;
 wire \requested_addr_latch[3] ;
 wire \requested_addr_latch[4] ;
 wire \requested_addr_latch[5] ;
 wire \requested_addr_latch[6] ;
 wire \requested_addr_latch[7] ;
 wire \requested_addr_latch[8] ;
 wire \requested_addr_latch[9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A4 (.I(net52),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__B2 (.I(_076_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__I (.I(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__B2 (.I(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__C1 (.I(net61),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__A4 (.I(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__115__A2 (.I(net37),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__116__A4 (.I(net53),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__118__B2 (.I(_083_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__I (.I(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__B2 (.I(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__C1 (.I(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__A4 (.I(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__A2 (.I(net38),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__A4 (.I(net54),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__B2 (.I(_090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__B2 (.I(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__C1 (.I(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__A4 (.I(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__A2 (.I(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__A4 (.I(net55),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__B2 (.I(_097_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__B2 (.I(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__C1 (.I(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__A4 (.I(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__A3 (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__A2 (.I(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__B (.I(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__A4 (.I(net56),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A1 (.I(_098_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A2 (.I(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__B2 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__A1 (.I(net74),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__A1 (.I(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__I (.I(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__I (.I(\requested_addr_latch[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__I (.I(\requested_addr_latch[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__I (.I(\requested_addr_latch[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I (.I(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__I (.I(\requested_addr_latch[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__I (.I(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__A4 (.I(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__A1 (.I(\requested_addr_latch[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__A2 (.I(\requested_addr_latch[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__I (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A2 (.I(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I (.I(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__A2 (.I(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__A4 (.I(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__A2 (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__I (.I(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__B2 (.I(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__C1 (.I(net57),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__A4 (.I(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__A4 (.I(net49),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__I (.I(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__B2 (.I(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__C1 (.I(net58),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__A4 (.I(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__A4 (.I(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I (.I(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__B2 (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__C1 (.I(net59),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__A4 (.I(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A2 (.I(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__A4 (.I(net51),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__B2 (.I(_059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__I (.I(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__I (.I(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__B2 (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__C1 (.I(net60),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__A4 (.I(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I (.I(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__I (.I(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__A2 (.I(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__D (.I(net75),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__D (.I(net82),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__D (.I(net83),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__CLK (.I(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__D (.I(net84),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__CLK (.I(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__D (.I(net85),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__CLK (.I(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__D (.I(net86),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__CLK (.I(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__D (.I(net87),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__CLK (.I(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__D (.I(net88),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__CLK (.I(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__D (.I(net89),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__CLK (.I(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__D (.I(net90),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__D (.I(net76),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__D (.I(net77),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__CLK (.I(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__I (.I(net84),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__I (.I(net85),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__I (.I(net86),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__I (.I(net87),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I (.I(net88),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__I (.I(net89),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__I (.I(net90),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__I (.I(net76),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__I (.I(net77),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__I (.I(net91),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I (.I(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__I (.I(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__I (.I(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__I (.I(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I (.I(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__I (.I(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I (.I(net72),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__I (.I(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(Q1[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(Q1[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(Q1[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(Q1[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(Q1[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(Q1[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(Q1[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(Q2[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(Q2[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(Q2[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(Q0[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(Q2[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(Q2[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(Q2[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(Q2[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(Q2[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(Q3[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(Q3[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(Q3[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(Q3[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(Q3[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(Q0[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(Q3[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(Q3[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(Q3[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(Q4[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(Q4[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(Q4[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(Q4[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(Q4[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(Q4[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(Q4[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(Q0[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(Q4[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(Q5[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(Q5[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(Q5[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(Q5[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(Q5[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(Q5[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(Q5[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(Q5[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(Q6[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(Q0[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(Q6[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(Q6[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(Q6[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(Q6[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(Q6[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(Q6[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(Q6[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(Q7[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(Q7[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(Q7[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(Q0[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(Q7[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(Q7[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(Q7[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(Q7[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(Q7[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(WEb_ram),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(bus_in[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(bus_in[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(bus_in[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(bus_in[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(Q0[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(bus_in[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(bus_in[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(bus_in[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(bus_in[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(ram_enabled),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(requested_addr[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(requested_addr[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(requested_addr[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(requested_addr[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(requested_addr[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(Q0[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(requested_addr[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(requested_addr[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(requested_addr[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(requested_addr[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(requested_addr[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(requested_addr[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(requested_addr[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(requested_addr[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(requested_addr[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(requested_addr[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(Q0[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(requested_addr[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(rst),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(Q1[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1002 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1019 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1022 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1026 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1035 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1051 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1062 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1070 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1074 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1083 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1090 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1098 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1491 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1515 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1532 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1563 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1566 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1574 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1578 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1587 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1595 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1600 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1602 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1611 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1650 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1659 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1665 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1668 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1672 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1674 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1691 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1695 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1697 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1708 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1716 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1720 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1722 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1733 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1736 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1744 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1757 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1765 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1770 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1797 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1799 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1812 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1818 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1829 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1833 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1835 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1838 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1853 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1861 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1865 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1867 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1880 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1888 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1890 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1901 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1903 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1914 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1925 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1933 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_575 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_610 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_618 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_674 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_678 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_716 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_743 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_750 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_754 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_784 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_786 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_795 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_811 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_813 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_824 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_832 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_834 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_843 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_847 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_849 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_852 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_856 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_858 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_867 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_875 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_879 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_881 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_900 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_904 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_915 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_917 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_920 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_928 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_930 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_939 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_949 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_954 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_956 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_963 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_979 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_983 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_994 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1433 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1455 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1491 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1468 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1456 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_455 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_596 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_623 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_668 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_695 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_710 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_716 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_732 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_740 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_767 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_769 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_776 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_780 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_784 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_832 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1007 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1033 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1035 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1044 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1048 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1064 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1068 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1077 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1479 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_520 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_529 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_560 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_584 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_599 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_608 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_823 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_827 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_843 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_855 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_864 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_868 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_872 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_874 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_885 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_897 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_901 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_917 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_925 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_955 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_959 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_975 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_979 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_995 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1068 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_858 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_860 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_890 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_894 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_898 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1002 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1010 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1014 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1033 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1037 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1069 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1073 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_815 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_819 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_849 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_853 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_873 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_893 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_923 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_931 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_939 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_943 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_963 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_994 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_998 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1033 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1037 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1045 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_928 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_963 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_967 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_971 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_998 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1032 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1036 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1044 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1048 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1468 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1433 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1463 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1258 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_660 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_689 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_693 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_697 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1010 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1022 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1029 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1045 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1049 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1051 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1056 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1058 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1065 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1085 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1090 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1092 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1520 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1538 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1554 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1572 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1588 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1622 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1634 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1657 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1668 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1670 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1695 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1699 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1704 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1715 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1733 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1736 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1740 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1751 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1767 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1770 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1774 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1776 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1795 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1799 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1804 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1812 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1823 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1831 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1835 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1838 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1846 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1848 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1859 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1867 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1869 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1872 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1880 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1884 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1901 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1903 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1914 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1918 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1920 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_509 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_550 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_584 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_618 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_652 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_668 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_690 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_694 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_705 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_713 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_716 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_732 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_741 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_745 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_747 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_750 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_768 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_777 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_784 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_800 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_804 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_813 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_815 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_818 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_834 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_838 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_840 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_849 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_852 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_868 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_876 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_880 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_908 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_926 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_942 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_960 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_994 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1491 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1392 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1017 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1081 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1087 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1717 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1781 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1787 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1851 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1857 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1921 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1927 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1935 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1937 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_731 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_737 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_807 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_871 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_947 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1046 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1052 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1458 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1752 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1816 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1822 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1886 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1892 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1924 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1932 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1936 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_702 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_766 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_772 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_912 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_982 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _106_ (.I(_004_),
    .Z(_073_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _107_ (.I(_025_),
    .Z(_074_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _108_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net52),
    .ZN(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _109_ (.A1(_068_),
    .A2(_070_),
    .A3(_072_),
    .A4(_075_),
    .Z(_076_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _110_ (.A1(_060_),
    .A2(_061_),
    .B1(_065_),
    .B2(_076_),
    .ZN(net121),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _111_ (.I(net5),
    .ZN(_077_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _112_ (.A1(net21),
    .A2(_062_),
    .B1(_063_),
    .B2(net45),
    .C1(net61),
    .C2(_064_),
    .ZN(_078_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _113_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net13),
    .ZN(_079_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _114_ (.A1(_053_),
    .A2(net29),
    .A3(_069_),
    .ZN(_080_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _115_ (.A1(_055_),
    .A2(net37),
    .B(_071_),
    .ZN(_081_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _116_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net53),
    .ZN(_082_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _117_ (.A1(_079_),
    .A2(_080_),
    .A3(_081_),
    .A4(_082_),
    .Z(_083_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _118_ (.A1(_077_),
    .A2(_061_),
    .B1(_078_),
    .B2(_083_),
    .ZN(net122),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _119_ (.I(net6),
    .ZN(_084_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _120_ (.A1(net22),
    .A2(_062_),
    .B1(_063_),
    .B2(net46),
    .C1(net62),
    .C2(_064_),
    .ZN(_085_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _121_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net14),
    .ZN(_086_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _122_ (.A1(_053_),
    .A2(net30),
    .A3(_069_),
    .ZN(_087_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _123_ (.A1(_055_),
    .A2(net38),
    .B(_071_),
    .ZN(_088_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _124_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net54),
    .ZN(_089_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _125_ (.A1(_086_),
    .A2(_087_),
    .A3(_088_),
    .A4(_089_),
    .Z(_090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _126_ (.A1(_084_),
    .A2(_061_),
    .B1(_085_),
    .B2(_090_),
    .ZN(net123),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _127_ (.I(net7),
    .ZN(_091_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _128_ (.A1(net23),
    .A2(_062_),
    .B1(_063_),
    .B2(net47),
    .C1(net63),
    .C2(_064_),
    .ZN(_092_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _129_ (.A1(_066_),
    .A2(_067_),
    .A3(_015_),
    .A4(net15),
    .ZN(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _130_ (.A1(_038_),
    .A2(net31),
    .A3(_069_),
    .ZN(_094_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _131_ (.A1(_035_),
    .A2(net39),
    .B(_071_),
    .ZN(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _132_ (.A1(_073_),
    .A2(_074_),
    .A3(_008_),
    .A4(net55),
    .ZN(_096_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _133_ (.A1(_093_),
    .A2(_094_),
    .A3(_095_),
    .A4(_096_),
    .Z(_097_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _134_ (.A1(_091_),
    .A2(_061_),
    .B1(_092_),
    .B2(_097_),
    .ZN(net124),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _135_ (.I(net8),
    .ZN(_098_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _136_ (.A1(net24),
    .A2(_018_),
    .B1(_026_),
    .B2(net48),
    .C1(net64),
    .C2(_030_),
    .ZN(_099_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _137_ (.A1(_011_),
    .A2(_006_),
    .A3(_015_),
    .A4(net16),
    .ZN(_100_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _138_ (.A1(_038_),
    .A2(net32),
    .A3(_020_),
    .ZN(_101_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _139_ (.A1(_035_),
    .A2(net40),
    .B(_023_),
    .ZN(_102_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _140_ (.A1(_004_),
    .A2(_025_),
    .A3(_008_),
    .A4(net56),
    .ZN(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _141_ (.A1(_100_),
    .A2(_101_),
    .A3(_102_),
    .A4(_103_),
    .Z(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _142_ (.A1(_098_),
    .A2(_009_),
    .B1(_099_),
    .B2(_104_),
    .ZN(net125),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _143_ (.A1(\requested_addr_latch[14] ),
    .A2(\requested_addr_latch[12] ),
    .A3(\requested_addr_latch[13] ),
    .ZN(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _144_ (.A1(net74),
    .A2(_105_),
    .ZN(_000_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _145_ (.A1(net65),
    .A2(\requested_addr_latch[15] ),
    .A3(_000_),
    .ZN(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _146_ (.I(_001_),
    .Z(_002_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _147_ (.I(\requested_addr_latch[1] ),
    .Z(_003_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _148_ (.I(_003_),
    .Z(_004_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _149_ (.I(\requested_addr_latch[0] ),
    .Z(_005_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _150_ (.I(_005_),
    .Z(_006_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _151_ (.I(\requested_addr_latch[2] ),
    .Z(_007_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _152_ (.I(_007_),
    .Z(_008_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _153_ (.A1(_004_),
    .A2(_006_),
    .A3(_008_),
    .ZN(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _154_ (.I(_009_),
    .Z(_010_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _155_ (.A1(_002_),
    .A2(_010_),
    .ZN(net110),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _156_ (.I(_003_),
    .ZN(_011_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _157_ (.I(_011_),
    .Z(_012_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _158_ (.I(_006_),
    .Z(_013_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _159_ (.I(\requested_addr_latch[2] ),
    .ZN(_014_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _160_ (.I(_014_),
    .Z(_015_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _161_ (.I(_015_),
    .Z(_016_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _162_ (.I(_001_),
    .Z(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _163_ (.A1(_012_),
    .A2(_013_),
    .A3(_016_),
    .A4(_017_),
    .ZN(net111),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _164_ (.A1(_011_),
    .A2(_005_),
    .A3(_007_),
    .ZN(_018_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _165_ (.I(_018_),
    .Z(_019_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _166_ (.A1(_002_),
    .A2(_019_),
    .ZN(net112),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _167_ (.A1(\requested_addr_latch[1] ),
    .A2(\requested_addr_latch[0] ),
    .Z(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _168_ (.I(_020_),
    .Z(_021_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _169_ (.A1(_016_),
    .A2(_017_),
    .A3(_021_),
    .ZN(net113),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _170_ (.I(_008_),
    .Z(_022_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _171_ (.A1(_003_),
    .A2(_005_),
    .ZN(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _172_ (.I(_023_),
    .Z(_024_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _173_ (.A1(_022_),
    .A2(_017_),
    .A3(_024_),
    .ZN(net114),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _174_ (.I(_005_),
    .ZN(_025_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _175_ (.A1(_003_),
    .A2(_025_),
    .A3(_014_),
    .ZN(_026_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _176_ (.I(_026_),
    .Z(_027_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _177_ (.A1(_002_),
    .A2(_027_),
    .ZN(net115),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _178_ (.I(_004_),
    .Z(_028_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _179_ (.I(_025_),
    .Z(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _180_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(_017_),
    .ZN(net116),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _181_ (.A1(_007_),
    .A2(_020_),
    .Z(_030_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _182_ (.I(_030_),
    .Z(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _183_ (.A1(_002_),
    .A2(_031_),
    .ZN(net117),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _184_ (.I(net1),
    .ZN(_032_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _185_ (.A1(net17),
    .A2(_019_),
    .B1(_027_),
    .B2(net41),
    .C1(net57),
    .C2(_031_),
    .ZN(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _186_ (.I(_014_),
    .Z(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _187_ (.I(_034_),
    .Z(_035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _188_ (.A1(_012_),
    .A2(_013_),
    .A3(_035_),
    .A4(net9),
    .ZN(_036_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _189_ (.A1(_016_),
    .A2(net25),
    .A3(_021_),
    .ZN(_037_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _190_ (.I(_034_),
    .Z(_038_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _191_ (.A1(_038_),
    .A2(net33),
    .B(_024_),
    .ZN(_039_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _192_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(net49),
    .ZN(_040_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _193_ (.A1(_036_),
    .A2(_037_),
    .A3(_039_),
    .A4(_040_),
    .Z(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _194_ (.A1(_032_),
    .A2(_010_),
    .B1(_033_),
    .B2(_041_),
    .ZN(net118),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _195_ (.I(net2),
    .ZN(_042_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _196_ (.A1(net18),
    .A2(_019_),
    .B1(_027_),
    .B2(net42),
    .C1(net58),
    .C2(_031_),
    .ZN(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _197_ (.A1(_012_),
    .A2(_013_),
    .A3(_035_),
    .A4(net10),
    .ZN(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _198_ (.A1(_016_),
    .A2(net26),
    .A3(_021_),
    .ZN(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _199_ (.A1(_038_),
    .A2(net34),
    .B(_024_),
    .ZN(_046_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _200_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(net50),
    .ZN(_047_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _201_ (.A1(_044_),
    .A2(_045_),
    .A3(_046_),
    .A4(_047_),
    .Z(_048_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _202_ (.A1(_042_),
    .A2(_010_),
    .B1(_043_),
    .B2(_048_),
    .ZN(net119),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _203_ (.I(net3),
    .ZN(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _204_ (.A1(net19),
    .A2(_019_),
    .B1(_027_),
    .B2(net43),
    .C1(net59),
    .C2(_031_),
    .ZN(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _205_ (.I(_034_),
    .Z(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _206_ (.A1(_012_),
    .A2(_013_),
    .A3(_051_),
    .A4(net11),
    .ZN(_052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _207_ (.I(_015_),
    .Z(_053_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _208_ (.A1(_053_),
    .A2(net27),
    .A3(_021_),
    .ZN(_054_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _209_ (.I(_034_),
    .Z(_055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _210_ (.A1(_055_),
    .A2(net35),
    .B(_024_),
    .ZN(_056_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _211_ (.I(_007_),
    .Z(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _212_ (.A1(_028_),
    .A2(_029_),
    .A3(_057_),
    .A4(net51),
    .ZN(_058_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _213_ (.A1(_052_),
    .A2(_054_),
    .A3(_056_),
    .A4(_058_),
    .Z(_059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _214_ (.A1(_049_),
    .A2(_010_),
    .B1(_050_),
    .B2(_059_),
    .ZN(net120),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _215_ (.I(net4),
    .ZN(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _216_ (.I(_009_),
    .Z(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _217_ (.I(_018_),
    .Z(_062_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _218_ (.I(_026_),
    .Z(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _219_ (.I(_030_),
    .Z(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _220_ (.A1(net20),
    .A2(_062_),
    .B1(_063_),
    .B2(net44),
    .C1(net60),
    .C2(_064_),
    .ZN(_065_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _221_ (.I(_011_),
    .Z(_066_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _222_ (.I(_006_),
    .Z(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _223_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net12),
    .ZN(_068_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _224_ (.I(_020_),
    .Z(_069_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _225_ (.A1(_053_),
    .A2(net28),
    .A3(_069_),
    .ZN(_070_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _226_ (.I(_023_),
    .Z(_071_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _227_ (.A1(_055_),
    .A2(net36),
    .B(_071_),
    .ZN(_072_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _228_ (.D(net75),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _229_ (.D(net82),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _230_ (.D(net83),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _231_ (.D(net84),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _232_ (.D(net85),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _233_ (.D(net86),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _234_ (.D(net87),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _235_ (.D(net88),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _236_ (.D(net89),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[8] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _237_ (.D(net90),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\requested_addr_latch[9] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _238_ (.D(net76),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[10] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _239_ (.D(net77),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[11] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _240_ (.D(net78),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[12] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _241_ (.D(net79),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[13] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _242_ (.D(net80),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[14] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _243_ (.D(net81),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\requested_addr_latch[15] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _252_ (.I(net84),
    .Z(net92),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _253_ (.I(net85),
    .Z(net93),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _254_ (.I(net86),
    .Z(net94),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _255_ (.I(net87),
    .Z(net95),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _256_ (.I(net88),
    .Z(net96),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _257_ (.I(net89),
    .Z(net97),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _258_ (.I(net90),
    .Z(net98),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _259_ (.I(net76),
    .Z(net99),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _260_ (.I(net77),
    .Z(net100),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _261_ (.I(net91),
    .Z(net101),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _262_ (.I(net66),
    .Z(net102),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _263_ (.I(net67),
    .Z(net103),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _264_ (.I(net68),
    .Z(net104),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _265_ (.I(net69),
    .Z(net105),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _266_ (.I(net70),
    .Z(net106),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _267_ (.I(net71),
    .Z(net107),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _268_ (.I(net72),
    .Z(net108),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _269_ (.I(net73),
    .Z(net109),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_0__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_1__leaf_wb_clk_i),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(Q0[0]),
    .Z(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(Q1[1]),
    .Z(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(Q1[2]),
    .Z(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(Q1[3]),
    .Z(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(Q1[4]),
    .Z(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(Q1[5]),
    .Z(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(Q1[6]),
    .Z(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(Q1[7]),
    .Z(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(Q2[0]),
    .Z(net17),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(Q2[1]),
    .Z(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(Q2[2]),
    .Z(net19),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(Q0[1]),
    .Z(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(Q2[3]),
    .Z(net20),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(Q2[4]),
    .Z(net21),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(Q2[5]),
    .Z(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(Q2[6]),
    .Z(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(Q2[7]),
    .Z(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(Q3[0]),
    .Z(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(Q3[1]),
    .Z(net26),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(Q3[2]),
    .Z(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(Q3[3]),
    .Z(net28),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(Q3[4]),
    .Z(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(Q0[2]),
    .Z(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(Q3[5]),
    .Z(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(Q3[6]),
    .Z(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(Q3[7]),
    .Z(net32),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(Q4[0]),
    .Z(net33),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(Q4[1]),
    .Z(net34),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(Q4[2]),
    .Z(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(Q4[3]),
    .Z(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(Q4[4]),
    .Z(net37),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(Q4[5]),
    .Z(net38),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(Q4[6]),
    .Z(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(Q0[3]),
    .Z(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(Q4[7]),
    .Z(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input41 (.I(Q5[0]),
    .Z(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input42 (.I(Q5[1]),
    .Z(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(Q5[2]),
    .Z(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input44 (.I(Q5[3]),
    .Z(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(Q5[4]),
    .Z(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(Q5[5]),
    .Z(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(Q5[6]),
    .Z(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(Q5[7]),
    .Z(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(Q6[0]),
    .Z(net49),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(Q0[4]),
    .Z(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(Q6[1]),
    .Z(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input51 (.I(Q6[2]),
    .Z(net51),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(Q6[3]),
    .Z(net52),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input53 (.I(Q6[4]),
    .Z(net53),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input54 (.I(Q6[5]),
    .Z(net54),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input55 (.I(Q6[6]),
    .Z(net55),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input56 (.I(Q6[7]),
    .Z(net56),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input57 (.I(Q7[0]),
    .Z(net57),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input58 (.I(Q7[1]),
    .Z(net58),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input59 (.I(Q7[2]),
    .Z(net59),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(Q0[5]),
    .Z(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input60 (.I(Q7[3]),
    .Z(net60),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input61 (.I(Q7[4]),
    .Z(net61),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input62 (.I(Q7[5]),
    .Z(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input63 (.I(Q7[6]),
    .Z(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input64 (.I(Q7[7]),
    .Z(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input65 (.I(WEb_ram),
    .Z(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input66 (.I(bus_in[0]),
    .Z(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input67 (.I(bus_in[1]),
    .Z(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input68 (.I(bus_in[2]),
    .Z(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input69 (.I(bus_in[3]),
    .Z(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(Q0[6]),
    .Z(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input70 (.I(bus_in[4]),
    .Z(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input71 (.I(bus_in[5]),
    .Z(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input72 (.I(bus_in[6]),
    .Z(net72),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input73 (.I(bus_in[7]),
    .Z(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input74 (.I(ram_enabled),
    .Z(net74),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input75 (.I(requested_addr[0]),
    .Z(net75),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input76 (.I(requested_addr[10]),
    .Z(net76),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input77 (.I(requested_addr[11]),
    .Z(net77),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(requested_addr[12]),
    .Z(net78),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(requested_addr[13]),
    .Z(net79),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(Q0[7]),
    .Z(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(requested_addr[14]),
    .Z(net80),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(requested_addr[15]),
    .Z(net81),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input82 (.I(requested_addr[1]),
    .Z(net82),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input83 (.I(requested_addr[2]),
    .Z(net83),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input84 (.I(requested_addr[3]),
    .Z(net84),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input85 (.I(requested_addr[4]),
    .Z(net85),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input86 (.I(requested_addr[5]),
    .Z(net86),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input87 (.I(requested_addr[6]),
    .Z(net87),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input88 (.I(requested_addr[7]),
    .Z(net88),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input89 (.I(requested_addr[8]),
    .Z(net89),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(Q1[0]),
    .Z(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input90 (.I(requested_addr[9]),
    .Z(net90),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input91 (.I(rst),
    .Z(net91),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output100 (.I(net100),
    .Z(A_all[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output101 (.I(net101),
    .Z(CEN_all),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output102 (.I(net102),
    .Z(D_all[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output103 (.I(net103),
    .Z(D_all[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output104 (.I(net104),
    .Z(D_all[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output105 (.I(net105),
    .Z(D_all[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(D_all[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(D_all[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(D_all[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(D_all[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(GWEN_0),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(GWEN_1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(GWEN_2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(GWEN_3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(GWEN_4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(GWEN_5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(GWEN_6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(GWEN_7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(bus_out[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(bus_out[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(bus_out[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(bus_out[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(bus_out[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(bus_out[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(bus_out[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(bus_out[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output92 (.I(net92),
    .Z(A_all[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output93 (.I(net93),
    .Z(A_all[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output94 (.I(net94),
    .Z(A_all[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output95 (.I(net95),
    .Z(A_all[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output96 (.I(net96),
    .Z(A_all[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output97 (.I(net97),
    .Z(A_all[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output98 (.I(net98),
    .Z(A_all[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output99 (.I(net99),
    .Z(A_all[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_126 (.ZN(net126),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_127 (.ZN(net127),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_128 (.ZN(net128),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_129 (.ZN(net129),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_130 (.ZN(net130),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_131 (.ZN(net131),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_132 (.ZN(net132),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_133 (.ZN(net133),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 assign WEN_all[0] = net126;
 assign WEN_all[1] = net127;
 assign WEN_all[2] = net128;
 assign WEN_all[3] = net129;
 assign WEN_all[4] = net130;
 assign WEN_all[5] = net131;
 assign WEN_all[6] = net132;
 assign WEN_all[7] = net133;
endmodule
