magic
tech gf180mcuD
magscale 1 10
timestamp 1700263339
<< metal1 >>
rect 38770 56590 38782 56642
rect 38834 56639 38846 56642
rect 39330 56639 39342 56642
rect 38834 56593 39342 56639
rect 38834 56590 38846 56593
rect 39330 56590 39342 56593
rect 39394 56639 39406 56642
rect 40114 56639 40126 56642
rect 39394 56593 40126 56639
rect 39394 56590 39406 56593
rect 40114 56590 40126 56593
rect 40178 56590 40190 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 5070 56306 5122 56318
rect 5070 56242 5122 56254
rect 7422 56306 7474 56318
rect 7422 56242 7474 56254
rect 7646 56306 7698 56318
rect 7646 56242 7698 56254
rect 9662 56306 9714 56318
rect 9662 56242 9714 56254
rect 9886 56306 9938 56318
rect 9886 56242 9938 56254
rect 11902 56306 11954 56318
rect 11902 56242 11954 56254
rect 12126 56306 12178 56318
rect 12126 56242 12178 56254
rect 14142 56306 14194 56318
rect 14142 56242 14194 56254
rect 16494 56306 16546 56318
rect 16494 56242 16546 56254
rect 16942 56306 16994 56318
rect 16942 56242 16994 56254
rect 18622 56306 18674 56318
rect 18622 56242 18674 56254
rect 18846 56306 18898 56318
rect 18846 56242 18898 56254
rect 20302 56306 20354 56318
rect 20302 56242 20354 56254
rect 23102 56306 23154 56318
rect 23102 56242 23154 56254
rect 25342 56306 25394 56318
rect 25342 56242 25394 56254
rect 29822 56306 29874 56318
rect 29822 56242 29874 56254
rect 31726 56306 31778 56318
rect 31726 56242 31778 56254
rect 34302 56306 34354 56318
rect 34302 56242 34354 56254
rect 36542 56306 36594 56318
rect 36542 56242 36594 56254
rect 39342 56306 39394 56318
rect 39342 56242 39394 56254
rect 41470 56306 41522 56318
rect 41470 56242 41522 56254
rect 44606 56306 44658 56318
rect 44606 56242 44658 56254
rect 48974 56306 49026 56318
rect 48974 56242 49026 56254
rect 52222 56306 52274 56318
rect 52222 56242 52274 56254
rect 56030 56306 56082 56318
rect 56030 56242 56082 56254
rect 2046 56194 2098 56206
rect 2046 56130 2098 56142
rect 2382 56194 2434 56206
rect 2382 56130 2434 56142
rect 5518 56194 5570 56206
rect 5518 56130 5570 56142
rect 5854 56194 5906 56206
rect 14366 56194 14418 56206
rect 21086 56194 21138 56206
rect 7970 56142 7982 56194
rect 8034 56142 8046 56194
rect 10210 56142 10222 56194
rect 10274 56142 10286 56194
rect 12450 56142 12462 56194
rect 12514 56142 12526 56194
rect 17266 56142 17278 56194
rect 17330 56142 17342 56194
rect 19170 56142 19182 56194
rect 19234 56142 19246 56194
rect 5854 56130 5906 56142
rect 14366 56130 14418 56142
rect 21086 56130 21138 56142
rect 21422 56194 21474 56206
rect 21422 56130 21474 56142
rect 23326 56194 23378 56206
rect 23326 56130 23378 56142
rect 25566 56194 25618 56206
rect 25566 56130 25618 56142
rect 28366 56194 28418 56206
rect 28366 56130 28418 56142
rect 30046 56194 30098 56206
rect 30046 56130 30098 56142
rect 32286 56194 32338 56206
rect 32286 56130 32338 56142
rect 32622 56194 32674 56206
rect 32622 56130 32674 56142
rect 34526 56194 34578 56206
rect 34526 56130 34578 56142
rect 34862 56194 34914 56206
rect 34862 56130 34914 56142
rect 36766 56194 36818 56206
rect 36766 56130 36818 56142
rect 37102 56194 37154 56206
rect 37102 56130 37154 56142
rect 39790 56194 39842 56206
rect 39790 56130 39842 56142
rect 40126 56194 40178 56206
rect 40126 56130 40178 56142
rect 1710 56082 1762 56094
rect 47742 56082 47794 56094
rect 54574 56082 54626 56094
rect 2594 56030 2606 56082
rect 2658 56030 2670 56082
rect 14578 56030 14590 56082
rect 14642 56030 14654 56082
rect 23538 56030 23550 56082
rect 23602 56030 23614 56082
rect 25778 56030 25790 56082
rect 25842 56030 25854 56082
rect 28578 56030 28590 56082
rect 28642 56030 28654 56082
rect 30258 56030 30270 56082
rect 30322 56030 30334 56082
rect 40450 56030 40462 56082
rect 40514 56030 40526 56082
rect 43698 56030 43710 56082
rect 43762 56030 43774 56082
rect 47954 56030 47966 56082
rect 48018 56030 48030 56082
rect 51202 56030 51214 56082
rect 51266 56030 51278 56082
rect 55010 56030 55022 56082
rect 55074 56030 55086 56082
rect 1710 56018 1762 56030
rect 47742 56018 47794 56030
rect 54574 56018 54626 56030
rect 3166 55970 3218 55982
rect 3166 55906 3218 55918
rect 27918 55970 27970 55982
rect 27918 55906 27970 55918
rect 38894 55970 38946 55982
rect 38894 55906 38946 55918
rect 27570 55806 27582 55858
rect 27634 55855 27646 55858
rect 27906 55855 27918 55858
rect 27634 55809 27918 55855
rect 27634 55806 27646 55809
rect 27906 55806 27918 55809
rect 27970 55806 27982 55858
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 2158 55410 2210 55422
rect 39118 55410 39170 55422
rect 46734 55410 46786 55422
rect 16370 55358 16382 55410
rect 16434 55358 16446 55410
rect 20514 55358 20526 55410
rect 20578 55358 20590 55410
rect 32050 55358 32062 55410
rect 32114 55358 32126 55410
rect 36418 55358 36430 55410
rect 36482 55358 36494 55410
rect 43138 55358 43150 55410
rect 43202 55358 43214 55410
rect 2158 55346 2210 55358
rect 39118 55346 39170 55358
rect 46734 55346 46786 55358
rect 53678 55410 53730 55422
rect 56690 55358 56702 55410
rect 56754 55358 56766 55410
rect 53678 55346 53730 55358
rect 16830 55298 16882 55310
rect 21422 55298 21474 55310
rect 13570 55246 13582 55298
rect 13634 55246 13646 55298
rect 17714 55246 17726 55298
rect 17778 55246 17790 55298
rect 16830 55234 16882 55246
rect 21422 55234 21474 55246
rect 22990 55298 23042 55310
rect 22990 55234 23042 55246
rect 25454 55298 25506 55310
rect 25454 55234 25506 55246
rect 27694 55298 27746 55310
rect 29250 55246 29262 55298
rect 29314 55246 29326 55298
rect 32610 55246 32622 55298
rect 32674 55246 32686 55298
rect 33618 55246 33630 55298
rect 33682 55246 33694 55298
rect 37090 55246 37102 55298
rect 37154 55246 37166 55298
rect 38322 55246 38334 55298
rect 38386 55246 38398 55298
rect 40226 55246 40238 55298
rect 40290 55246 40302 55298
rect 45714 55246 45726 55298
rect 45778 55246 45790 55298
rect 52658 55246 52670 55298
rect 52722 55246 52734 55298
rect 55570 55246 55582 55298
rect 55634 55246 55646 55298
rect 27694 55234 27746 55246
rect 11790 55186 11842 55198
rect 14242 55134 14254 55186
rect 14306 55134 14318 55186
rect 18386 55134 18398 55186
rect 18450 55134 18462 55186
rect 29922 55134 29934 55186
rect 29986 55134 29998 55186
rect 34290 55134 34302 55186
rect 34354 55134 34366 55186
rect 37314 55134 37326 55186
rect 37378 55134 37390 55186
rect 41010 55134 41022 55186
rect 41074 55134 41086 55186
rect 11790 55122 11842 55134
rect 11902 55074 11954 55086
rect 11902 55010 11954 55022
rect 22878 55074 22930 55086
rect 22878 55010 22930 55022
rect 25342 55074 25394 55086
rect 25342 55010 25394 55022
rect 27582 55074 27634 55086
rect 27582 55010 27634 55022
rect 32622 55074 32674 55086
rect 32622 55010 32674 55022
rect 33182 55074 33234 55086
rect 33182 55010 33234 55022
rect 37774 55074 37826 55086
rect 39006 55074 39058 55086
rect 38098 55022 38110 55074
rect 38162 55022 38174 55074
rect 37774 55010 37826 55022
rect 39006 55010 39058 55022
rect 39902 55074 39954 55086
rect 39902 55010 39954 55022
rect 43598 55074 43650 55086
rect 43598 55010 43650 55022
rect 45390 55074 45442 55086
rect 45390 55010 45442 55022
rect 50878 55074 50930 55086
rect 50878 55010 50930 55022
rect 52110 55074 52162 55086
rect 52110 55010 52162 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 14702 54738 14754 54750
rect 14702 54674 14754 54686
rect 15822 54738 15874 54750
rect 15822 54674 15874 54686
rect 17614 54738 17666 54750
rect 17614 54674 17666 54686
rect 18510 54738 18562 54750
rect 18510 54674 18562 54686
rect 29486 54738 29538 54750
rect 29486 54674 29538 54686
rect 29934 54738 29986 54750
rect 29934 54674 29986 54686
rect 32510 54738 32562 54750
rect 32510 54674 32562 54686
rect 33966 54738 34018 54750
rect 33966 54674 34018 54686
rect 41022 54738 41074 54750
rect 41022 54674 41074 54686
rect 2046 54626 2098 54638
rect 15150 54626 15202 54638
rect 12786 54574 12798 54626
rect 12850 54574 12862 54626
rect 13122 54574 13134 54626
rect 13186 54574 13198 54626
rect 2046 54562 2098 54574
rect 15150 54562 15202 54574
rect 29150 54626 29202 54638
rect 29150 54562 29202 54574
rect 31838 54626 31890 54638
rect 36206 54626 36258 54638
rect 33394 54574 33406 54626
rect 33458 54574 33470 54626
rect 31838 54562 31890 54574
rect 36206 54562 36258 54574
rect 38894 54626 38946 54638
rect 38894 54562 38946 54574
rect 39566 54626 39618 54638
rect 39566 54562 39618 54574
rect 40910 54626 40962 54638
rect 40910 54562 40962 54574
rect 1710 54514 1762 54526
rect 1710 54450 1762 54462
rect 12462 54514 12514 54526
rect 14590 54514 14642 54526
rect 13682 54462 13694 54514
rect 13746 54462 13758 54514
rect 12462 54450 12514 54462
rect 14590 54450 14642 54462
rect 14926 54514 14978 54526
rect 14926 54450 14978 54462
rect 15710 54514 15762 54526
rect 15710 54450 15762 54462
rect 15934 54514 15986 54526
rect 15934 54450 15986 54462
rect 16382 54514 16434 54526
rect 16382 54450 16434 54462
rect 17278 54514 17330 54526
rect 17278 54450 17330 54462
rect 17614 54514 17666 54526
rect 17614 54450 17666 54462
rect 17838 54514 17890 54526
rect 17838 54450 17890 54462
rect 18286 54514 18338 54526
rect 18286 54450 18338 54462
rect 18398 54514 18450 54526
rect 28814 54514 28866 54526
rect 18834 54462 18846 54514
rect 18898 54462 18910 54514
rect 20962 54462 20974 54514
rect 21026 54462 21038 54514
rect 25218 54462 25230 54514
rect 25282 54462 25294 54514
rect 18398 54450 18450 54462
rect 28814 54450 28866 54462
rect 29822 54514 29874 54526
rect 33182 54514 33234 54526
rect 38222 54514 38274 54526
rect 30034 54462 30046 54514
rect 30098 54462 30110 54514
rect 30594 54462 30606 54514
rect 30658 54462 30670 54514
rect 33954 54462 33966 54514
rect 34018 54462 34030 54514
rect 34850 54462 34862 54514
rect 34914 54462 34926 54514
rect 29822 54450 29874 54462
rect 33182 54450 33234 54462
rect 38222 54450 38274 54462
rect 38558 54514 38610 54526
rect 38558 54450 38610 54462
rect 39230 54514 39282 54526
rect 41358 54514 41410 54526
rect 41122 54462 41134 54514
rect 41186 54462 41198 54514
rect 41458 54462 41470 54514
rect 41522 54462 41534 54514
rect 39230 54450 39282 54462
rect 41358 54450 41410 54462
rect 2494 54402 2546 54414
rect 36878 54402 36930 54414
rect 13794 54350 13806 54402
rect 13858 54350 13870 54402
rect 21746 54350 21758 54402
rect 21810 54350 21822 54402
rect 23874 54350 23886 54402
rect 23938 54350 23950 54402
rect 26002 54350 26014 54402
rect 26066 54350 26078 54402
rect 28130 54350 28142 54402
rect 28194 54350 28206 54402
rect 31714 54350 31726 54402
rect 31778 54350 31790 54402
rect 34738 54350 34750 54402
rect 34802 54350 34814 54402
rect 36082 54350 36094 54402
rect 36146 54350 36158 54402
rect 2494 54338 2546 54350
rect 36878 54338 36930 54350
rect 40350 54402 40402 54414
rect 40350 54338 40402 54350
rect 55246 54402 55298 54414
rect 55246 54338 55298 54350
rect 32062 54290 32114 54302
rect 30370 54238 30382 54290
rect 30434 54238 30446 54290
rect 32062 54226 32114 54238
rect 33630 54290 33682 54302
rect 33630 54226 33682 54238
rect 36430 54290 36482 54302
rect 36430 54226 36482 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 40910 53954 40962 53966
rect 40910 53890 40962 53902
rect 41246 53954 41298 53966
rect 41246 53890 41298 53902
rect 23662 53842 23714 53854
rect 23662 53778 23714 53790
rect 26350 53842 26402 53854
rect 26350 53778 26402 53790
rect 29262 53842 29314 53854
rect 29262 53778 29314 53790
rect 37662 53842 37714 53854
rect 37662 53778 37714 53790
rect 38894 53842 38946 53854
rect 42018 53790 42030 53842
rect 42082 53790 42094 53842
rect 38894 53778 38946 53790
rect 18174 53730 18226 53742
rect 16370 53678 16382 53730
rect 16434 53678 16446 53730
rect 18174 53666 18226 53678
rect 21982 53730 22034 53742
rect 21982 53666 22034 53678
rect 22430 53730 22482 53742
rect 22430 53666 22482 53678
rect 22654 53730 22706 53742
rect 22654 53666 22706 53678
rect 22878 53730 22930 53742
rect 22878 53666 22930 53678
rect 24446 53730 24498 53742
rect 24446 53666 24498 53678
rect 25118 53730 25170 53742
rect 33058 53678 33070 53730
rect 33122 53678 33134 53730
rect 38210 53678 38222 53730
rect 38274 53678 38286 53730
rect 41234 53678 41246 53730
rect 41298 53678 41310 53730
rect 25118 53666 25170 53678
rect 22318 53618 22370 53630
rect 16594 53566 16606 53618
rect 16658 53566 16670 53618
rect 22318 53554 22370 53566
rect 24894 53618 24946 53630
rect 24894 53554 24946 53566
rect 32622 53618 32674 53630
rect 32622 53554 32674 53566
rect 33294 53618 33346 53630
rect 33294 53554 33346 53566
rect 42366 53618 42418 53630
rect 42366 53554 42418 53566
rect 10446 53506 10498 53518
rect 10446 53442 10498 53454
rect 11566 53506 11618 53518
rect 11566 53442 11618 53454
rect 15374 53506 15426 53518
rect 15374 53442 15426 53454
rect 15934 53506 15986 53518
rect 15934 53442 15986 53454
rect 23550 53506 23602 53518
rect 23550 53442 23602 53454
rect 23774 53506 23826 53518
rect 23774 53442 23826 53454
rect 23998 53506 24050 53518
rect 23998 53442 24050 53454
rect 24782 53506 24834 53518
rect 24782 53442 24834 53454
rect 25566 53506 25618 53518
rect 25566 53442 25618 53454
rect 26238 53506 26290 53518
rect 26238 53442 26290 53454
rect 26462 53506 26514 53518
rect 26462 53442 26514 53454
rect 26686 53506 26738 53518
rect 42142 53506 42194 53518
rect 37986 53454 37998 53506
rect 38050 53454 38062 53506
rect 26686 53442 26738 53454
rect 42142 53442 42194 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 12798 53170 12850 53182
rect 12798 53106 12850 53118
rect 23438 53170 23490 53182
rect 23438 53106 23490 53118
rect 29150 53170 29202 53182
rect 29150 53106 29202 53118
rect 31950 53170 32002 53182
rect 31950 53106 32002 53118
rect 33854 53170 33906 53182
rect 41346 53118 41358 53170
rect 41410 53118 41422 53170
rect 33854 53106 33906 53118
rect 2046 53058 2098 53070
rect 9886 53058 9938 53070
rect 7970 53006 7982 53058
rect 8034 53006 8046 53058
rect 2046 52994 2098 53006
rect 9886 52994 9938 53006
rect 10670 53058 10722 53070
rect 10670 52994 10722 53006
rect 12014 53058 12066 53070
rect 12014 52994 12066 53006
rect 12350 53058 12402 53070
rect 12350 52994 12402 53006
rect 22766 53058 22818 53070
rect 29598 53058 29650 53070
rect 26674 53006 26686 53058
rect 26738 53006 26750 53058
rect 22766 52994 22818 53006
rect 29598 52994 29650 53006
rect 29934 53058 29986 53070
rect 32174 53058 32226 53070
rect 30146 53006 30158 53058
rect 30210 53006 30222 53058
rect 29934 52994 29986 53006
rect 32174 52994 32226 53006
rect 33070 53058 33122 53070
rect 33070 52994 33122 53006
rect 36430 53058 36482 53070
rect 36430 52994 36482 53006
rect 36542 53058 36594 53070
rect 36542 52994 36594 53006
rect 40910 53058 40962 53070
rect 42802 53006 42814 53058
rect 42866 53006 42878 53058
rect 40910 52994 40962 53006
rect 1710 52946 1762 52958
rect 10222 52946 10274 52958
rect 8754 52894 8766 52946
rect 8818 52894 8830 52946
rect 1710 52882 1762 52894
rect 10222 52882 10274 52894
rect 10558 52946 10610 52958
rect 10558 52882 10610 52894
rect 10894 52946 10946 52958
rect 17950 52946 18002 52958
rect 11330 52894 11342 52946
rect 11394 52894 11406 52946
rect 10894 52882 10946 52894
rect 17950 52882 18002 52894
rect 18398 52946 18450 52958
rect 18398 52882 18450 52894
rect 18510 52946 18562 52958
rect 18510 52882 18562 52894
rect 22318 52946 22370 52958
rect 22318 52882 22370 52894
rect 22990 52946 23042 52958
rect 22990 52882 23042 52894
rect 25454 52946 25506 52958
rect 25454 52882 25506 52894
rect 25902 52946 25954 52958
rect 25902 52882 25954 52894
rect 26126 52946 26178 52958
rect 26126 52882 26178 52894
rect 27022 52946 27074 52958
rect 27022 52882 27074 52894
rect 30382 52946 30434 52958
rect 30706 52894 30718 52946
rect 30770 52894 30782 52946
rect 33282 52894 33294 52946
rect 33346 52894 33358 52946
rect 33842 52894 33854 52946
rect 33906 52894 33918 52946
rect 36754 52894 36766 52946
rect 36818 52894 36830 52946
rect 41122 52894 41134 52946
rect 41186 52894 41198 52946
rect 41682 52894 41694 52946
rect 41746 52894 41758 52946
rect 42018 52894 42030 52946
rect 42082 52894 42094 52946
rect 30382 52882 30434 52894
rect 2494 52834 2546 52846
rect 15374 52834 15426 52846
rect 5842 52782 5854 52834
rect 5906 52782 5918 52834
rect 2494 52770 2546 52782
rect 15374 52770 15426 52782
rect 18174 52834 18226 52846
rect 18174 52770 18226 52782
rect 19070 52834 19122 52846
rect 19070 52770 19122 52782
rect 22542 52834 22594 52846
rect 22542 52770 22594 52782
rect 26014 52834 26066 52846
rect 26014 52770 26066 52782
rect 27470 52834 27522 52846
rect 27470 52770 27522 52782
rect 30046 52834 30098 52846
rect 36206 52834 36258 52846
rect 31826 52782 31838 52834
rect 31890 52782 31902 52834
rect 30046 52770 30098 52782
rect 36206 52770 36258 52782
rect 40350 52834 40402 52846
rect 44930 52782 44942 52834
rect 44994 52782 45006 52834
rect 40350 52770 40402 52782
rect 11006 52722 11058 52734
rect 29486 52722 29538 52734
rect 37214 52722 37266 52734
rect 2258 52670 2270 52722
rect 2322 52719 2334 52722
rect 2594 52719 2606 52722
rect 2322 52673 2606 52719
rect 2322 52670 2334 52673
rect 2594 52670 2606 52673
rect 2658 52670 2670 52722
rect 25106 52670 25118 52722
rect 25170 52719 25182 52722
rect 25330 52719 25342 52722
rect 25170 52673 25342 52719
rect 25170 52670 25182 52673
rect 25330 52670 25342 52673
rect 25394 52670 25406 52722
rect 33618 52670 33630 52722
rect 33682 52670 33694 52722
rect 41458 52670 41470 52722
rect 41522 52670 41534 52722
rect 11006 52658 11058 52670
rect 29486 52658 29538 52670
rect 37214 52658 37266 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 10446 52386 10498 52398
rect 11666 52334 11678 52386
rect 11730 52334 11742 52386
rect 10446 52322 10498 52334
rect 12798 52274 12850 52286
rect 12798 52210 12850 52222
rect 15598 52274 15650 52286
rect 32734 52274 32786 52286
rect 36990 52274 37042 52286
rect 17826 52222 17838 52274
rect 17890 52222 17902 52274
rect 19954 52222 19966 52274
rect 20018 52222 20030 52274
rect 22082 52222 22094 52274
rect 22146 52222 22158 52274
rect 30146 52222 30158 52274
rect 30210 52222 30222 52274
rect 32274 52222 32286 52274
rect 32338 52222 32350 52274
rect 34066 52222 34078 52274
rect 34130 52222 34142 52274
rect 36194 52222 36206 52274
rect 36258 52222 36270 52274
rect 15598 52210 15650 52222
rect 32734 52210 32786 52222
rect 36990 52210 37042 52222
rect 37102 52274 37154 52286
rect 41246 52274 41298 52286
rect 38658 52222 38670 52274
rect 38722 52222 38734 52274
rect 42578 52222 42590 52274
rect 42642 52222 42654 52274
rect 37102 52210 37154 52222
rect 41246 52210 41298 52222
rect 8990 52162 9042 52174
rect 8990 52098 9042 52110
rect 9998 52162 10050 52174
rect 9998 52098 10050 52110
rect 10334 52162 10386 52174
rect 11118 52162 11170 52174
rect 12350 52162 12402 52174
rect 10770 52110 10782 52162
rect 10834 52110 10846 52162
rect 11330 52110 11342 52162
rect 11394 52110 11406 52162
rect 11890 52110 11902 52162
rect 11954 52110 11966 52162
rect 10334 52098 10386 52110
rect 11118 52098 11170 52110
rect 12350 52098 12402 52110
rect 14590 52162 14642 52174
rect 14590 52098 14642 52110
rect 14814 52162 14866 52174
rect 14814 52098 14866 52110
rect 15150 52162 15202 52174
rect 15150 52098 15202 52110
rect 15710 52162 15762 52174
rect 27470 52162 27522 52174
rect 42478 52162 42530 52174
rect 16034 52110 16046 52162
rect 16098 52110 16110 52162
rect 20738 52110 20750 52162
rect 20802 52110 20814 52162
rect 27010 52110 27022 52162
rect 27074 52110 27086 52162
rect 29362 52110 29374 52162
rect 29426 52110 29438 52162
rect 33394 52110 33406 52162
rect 33458 52110 33470 52162
rect 37314 52110 37326 52162
rect 37378 52110 37390 52162
rect 38210 52110 38222 52162
rect 38274 52110 38286 52162
rect 40226 52110 40238 52162
rect 40290 52110 40302 52162
rect 42914 52110 42926 52162
rect 42978 52110 42990 52162
rect 15710 52098 15762 52110
rect 27470 52098 27522 52110
rect 42478 52098 42530 52110
rect 42142 52050 42194 52062
rect 39106 51998 39118 52050
rect 39170 51998 39182 52050
rect 42142 51986 42194 51998
rect 10110 51938 10162 51950
rect 10110 51874 10162 51886
rect 11902 51938 11954 51950
rect 11902 51874 11954 51886
rect 14702 51938 14754 51950
rect 14702 51874 14754 51886
rect 15486 51938 15538 51950
rect 15486 51874 15538 51886
rect 41694 51938 41746 51950
rect 41694 51874 41746 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 12014 51602 12066 51614
rect 23102 51602 23154 51614
rect 16482 51550 16494 51602
rect 16546 51550 16558 51602
rect 12014 51538 12066 51550
rect 23102 51538 23154 51550
rect 38894 51602 38946 51614
rect 38894 51538 38946 51550
rect 40126 51602 40178 51614
rect 40126 51538 40178 51550
rect 42254 51602 42306 51614
rect 42254 51538 42306 51550
rect 2046 51490 2098 51502
rect 2046 51426 2098 51438
rect 10670 51490 10722 51502
rect 39678 51490 39730 51502
rect 10882 51438 10894 51490
rect 10946 51438 10958 51490
rect 13906 51438 13918 51490
rect 13970 51438 13982 51490
rect 18722 51438 18734 51490
rect 18786 51438 18798 51490
rect 10670 51426 10722 51438
rect 39678 51426 39730 51438
rect 40350 51490 40402 51502
rect 40350 51426 40402 51438
rect 41022 51490 41074 51502
rect 41234 51438 41246 51490
rect 41298 51438 41310 51490
rect 41022 51426 41074 51438
rect 7646 51378 7698 51390
rect 1810 51326 1822 51378
rect 1874 51326 1886 51378
rect 4386 51326 4398 51378
rect 4450 51326 4462 51378
rect 7646 51314 7698 51326
rect 11118 51378 11170 51390
rect 16830 51378 16882 51390
rect 41470 51378 41522 51390
rect 11218 51326 11230 51378
rect 11282 51326 11294 51378
rect 13122 51326 13134 51378
rect 13186 51326 13198 51378
rect 22642 51326 22654 51378
rect 22706 51326 22718 51378
rect 25330 51326 25342 51378
rect 25394 51326 25406 51378
rect 39106 51326 39118 51378
rect 39170 51326 39182 51378
rect 39442 51326 39454 51378
rect 39506 51326 39518 51378
rect 41794 51326 41806 51378
rect 41858 51326 41870 51378
rect 11118 51314 11170 51326
rect 16830 51314 16882 51326
rect 41470 51314 41522 51326
rect 2494 51266 2546 51278
rect 10782 51266 10834 51278
rect 36430 51266 36482 51278
rect 5058 51214 5070 51266
rect 5122 51214 5134 51266
rect 7186 51214 7198 51266
rect 7250 51214 7262 51266
rect 16034 51214 16046 51266
rect 16098 51214 16110 51266
rect 26114 51214 26126 51266
rect 26178 51214 26190 51266
rect 28242 51214 28254 51266
rect 28306 51214 28318 51266
rect 2494 51202 2546 51214
rect 10782 51202 10834 51214
rect 36430 51202 36482 51214
rect 38558 51266 38610 51278
rect 38558 51202 38610 51214
rect 41134 51266 41186 51278
rect 42130 51214 42142 51266
rect 42194 51214 42206 51266
rect 41134 51202 41186 51214
rect 39230 51154 39282 51166
rect 39230 51090 39282 51102
rect 40014 51154 40066 51166
rect 40014 51090 40066 51102
rect 42478 51154 42530 51166
rect 42478 51090 42530 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 7310 50818 7362 50830
rect 7310 50754 7362 50766
rect 5070 50706 5122 50718
rect 1698 50654 1710 50706
rect 1762 50654 1774 50706
rect 3826 50654 3838 50706
rect 3890 50654 3902 50706
rect 5070 50642 5122 50654
rect 7086 50706 7138 50718
rect 7086 50642 7138 50654
rect 15934 50706 15986 50718
rect 15934 50642 15986 50654
rect 16494 50706 16546 50718
rect 16494 50642 16546 50654
rect 18286 50706 18338 50718
rect 26462 50706 26514 50718
rect 22082 50654 22094 50706
rect 22146 50654 22158 50706
rect 24210 50654 24222 50706
rect 24274 50654 24286 50706
rect 18286 50642 18338 50654
rect 26462 50642 26514 50654
rect 27358 50706 27410 50718
rect 27358 50642 27410 50654
rect 34638 50706 34690 50718
rect 37986 50654 37998 50706
rect 38050 50654 38062 50706
rect 40114 50654 40126 50706
rect 40178 50654 40190 50706
rect 44146 50654 44158 50706
rect 44210 50654 44222 50706
rect 34638 50642 34690 50654
rect 17390 50594 17442 50606
rect 4610 50542 4622 50594
rect 4674 50542 4686 50594
rect 17390 50530 17442 50542
rect 18174 50594 18226 50606
rect 18174 50530 18226 50542
rect 18846 50594 18898 50606
rect 25230 50594 25282 50606
rect 21410 50542 21422 50594
rect 21474 50542 21486 50594
rect 18846 50530 18898 50542
rect 25230 50530 25282 50542
rect 26238 50594 26290 50606
rect 26238 50530 26290 50542
rect 26686 50594 26738 50606
rect 26686 50530 26738 50542
rect 26798 50594 26850 50606
rect 26798 50530 26850 50542
rect 30270 50594 30322 50606
rect 36430 50594 36482 50606
rect 40910 50594 40962 50606
rect 35186 50542 35198 50594
rect 35250 50542 35262 50594
rect 37314 50542 37326 50594
rect 37378 50542 37390 50594
rect 41346 50542 41358 50594
rect 41410 50542 41422 50594
rect 30270 50530 30322 50542
rect 36430 50530 36482 50542
rect 40910 50530 40962 50542
rect 18398 50482 18450 50494
rect 17714 50430 17726 50482
rect 17778 50430 17790 50482
rect 18398 50418 18450 50430
rect 24782 50482 24834 50494
rect 25442 50430 25454 50482
rect 25506 50430 25518 50482
rect 42018 50430 42030 50482
rect 42082 50430 42094 50482
rect 24782 50418 24834 50430
rect 11902 50370 11954 50382
rect 7634 50318 7646 50370
rect 7698 50318 7710 50370
rect 11902 50306 11954 50318
rect 12574 50370 12626 50382
rect 12574 50306 12626 50318
rect 16046 50370 16098 50382
rect 16046 50306 16098 50318
rect 24558 50370 24610 50382
rect 24558 50306 24610 50318
rect 24670 50370 24722 50382
rect 24670 50306 24722 50318
rect 25790 50370 25842 50382
rect 32398 50370 32450 50382
rect 30594 50318 30606 50370
rect 30658 50318 30670 50370
rect 34962 50318 34974 50370
rect 35026 50318 35038 50370
rect 25790 50306 25842 50318
rect 32398 50306 32450 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 5070 50034 5122 50046
rect 5070 49970 5122 49982
rect 11342 50034 11394 50046
rect 11342 49970 11394 49982
rect 12014 50034 12066 50046
rect 12014 49970 12066 49982
rect 15262 50034 15314 50046
rect 33182 50034 33234 50046
rect 22418 49982 22430 50034
rect 22482 49982 22494 50034
rect 15262 49970 15314 49982
rect 33182 49970 33234 49982
rect 7198 49922 7250 49934
rect 3826 49870 3838 49922
rect 3890 49870 3902 49922
rect 7198 49858 7250 49870
rect 7534 49922 7586 49934
rect 25230 49922 25282 49934
rect 13122 49870 13134 49922
rect 13186 49870 13198 49922
rect 7534 49858 7586 49870
rect 25230 49858 25282 49870
rect 27582 49922 27634 49934
rect 27582 49858 27634 49870
rect 22094 49810 22146 49822
rect 4610 49758 4622 49810
rect 4674 49758 4686 49810
rect 6514 49758 6526 49810
rect 6578 49758 6590 49810
rect 8866 49758 8878 49810
rect 8930 49758 8942 49810
rect 10434 49758 10446 49810
rect 10498 49758 10510 49810
rect 11554 49758 11566 49810
rect 11618 49758 11630 49810
rect 12226 49758 12238 49810
rect 12290 49758 12302 49810
rect 12898 49758 12910 49810
rect 12962 49758 12974 49810
rect 32162 49758 32174 49810
rect 32226 49758 32238 49810
rect 37314 49758 37326 49810
rect 37378 49758 37390 49810
rect 22094 49746 22146 49758
rect 14926 49698 14978 49710
rect 1698 49646 1710 49698
rect 1762 49646 1774 49698
rect 6402 49646 6414 49698
rect 6466 49646 6478 49698
rect 6962 49646 6974 49698
rect 7026 49646 7038 49698
rect 7970 49646 7982 49698
rect 8034 49646 8046 49698
rect 8530 49646 8542 49698
rect 8594 49646 8606 49698
rect 10098 49646 10110 49698
rect 10162 49646 10174 49698
rect 14926 49634 14978 49646
rect 21758 49698 21810 49710
rect 21758 49634 21810 49646
rect 25790 49698 25842 49710
rect 37774 49698 37826 49710
rect 29250 49646 29262 49698
rect 29314 49646 29326 49698
rect 31378 49646 31390 49698
rect 31442 49646 31454 49698
rect 34402 49646 34414 49698
rect 34466 49646 34478 49698
rect 36530 49646 36542 49698
rect 36594 49646 36606 49698
rect 25790 49634 25842 49646
rect 37774 49634 37826 49646
rect 11230 49586 11282 49598
rect 11230 49522 11282 49534
rect 11902 49586 11954 49598
rect 11902 49522 11954 49534
rect 25342 49586 25394 49598
rect 25342 49522 25394 49534
rect 27694 49586 27746 49598
rect 27694 49522 27746 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 35858 49198 35870 49250
rect 35922 49247 35934 49250
rect 36530 49247 36542 49250
rect 35922 49201 36542 49247
rect 35922 49198 35934 49201
rect 36530 49198 36542 49201
rect 36594 49198 36606 49250
rect 10222 49138 10274 49150
rect 11902 49138 11954 49150
rect 6626 49086 6638 49138
rect 6690 49086 6702 49138
rect 11330 49086 11342 49138
rect 11394 49086 11406 49138
rect 10222 49074 10274 49086
rect 11902 49074 11954 49086
rect 12462 49138 12514 49150
rect 12462 49074 12514 49086
rect 14366 49138 14418 49150
rect 14366 49074 14418 49086
rect 15934 49138 15986 49150
rect 15934 49074 15986 49086
rect 19182 49138 19234 49150
rect 24558 49138 24610 49150
rect 35534 49138 35586 49150
rect 19954 49086 19966 49138
rect 20018 49086 20030 49138
rect 29586 49086 29598 49138
rect 29650 49086 29662 49138
rect 19182 49074 19234 49086
rect 24558 49074 24610 49086
rect 35534 49074 35586 49086
rect 38446 49138 38498 49150
rect 38446 49074 38498 49086
rect 7086 49026 7138 49038
rect 13918 49026 13970 49038
rect 11442 48974 11454 49026
rect 11506 48974 11518 49026
rect 7086 48962 7138 48974
rect 13918 48962 13970 48974
rect 14142 49026 14194 49038
rect 14142 48962 14194 48974
rect 15150 49026 15202 49038
rect 16494 49026 16546 49038
rect 15362 48974 15374 49026
rect 15426 48974 15438 49026
rect 15150 48962 15202 48974
rect 16494 48962 16546 48974
rect 17502 49026 17554 49038
rect 17502 48962 17554 48974
rect 18062 49026 18114 49038
rect 19406 49026 19458 49038
rect 19058 48974 19070 49026
rect 19122 48974 19134 49026
rect 18062 48962 18114 48974
rect 19406 48962 19458 48974
rect 20526 49026 20578 49038
rect 22094 49026 22146 49038
rect 21858 48974 21870 49026
rect 21922 48974 21934 49026
rect 20526 48962 20578 48974
rect 22094 48962 22146 48974
rect 22206 49026 22258 49038
rect 22206 48962 22258 48974
rect 24670 49026 24722 49038
rect 27918 49026 27970 49038
rect 32846 49026 32898 49038
rect 25666 48974 25678 49026
rect 25730 48974 25742 49026
rect 27122 48974 27134 49026
rect 27186 48974 27198 49026
rect 32498 48974 32510 49026
rect 32562 48974 32574 49026
rect 24670 48962 24722 48974
rect 27918 48962 27970 48974
rect 32846 48962 32898 48974
rect 34190 49026 34242 49038
rect 34190 48962 34242 48974
rect 34302 49026 34354 49038
rect 34302 48962 34354 48974
rect 35086 49026 35138 49038
rect 35086 48962 35138 48974
rect 35422 49026 35474 49038
rect 35422 48962 35474 48974
rect 1710 48914 1762 48926
rect 1710 48850 1762 48862
rect 11118 48914 11170 48926
rect 11118 48850 11170 48862
rect 16382 48914 16434 48926
rect 16382 48850 16434 48862
rect 17614 48914 17666 48926
rect 17614 48850 17666 48862
rect 17838 48914 17890 48926
rect 17838 48850 17890 48862
rect 19630 48914 19682 48926
rect 19630 48850 19682 48862
rect 19854 48914 19906 48926
rect 19854 48850 19906 48862
rect 20414 48914 20466 48926
rect 20414 48850 20466 48862
rect 22542 48914 22594 48926
rect 22542 48850 22594 48862
rect 22878 48914 22930 48926
rect 22878 48850 22930 48862
rect 22990 48914 23042 48926
rect 33070 48914 33122 48926
rect 25442 48862 25454 48914
rect 25506 48862 25518 48914
rect 27346 48862 27358 48914
rect 27410 48862 27422 48914
rect 31714 48862 31726 48914
rect 31778 48862 31790 48914
rect 22990 48850 23042 48862
rect 33070 48850 33122 48862
rect 35646 48914 35698 48926
rect 35646 48850 35698 48862
rect 2046 48802 2098 48814
rect 2046 48738 2098 48750
rect 2494 48802 2546 48814
rect 2494 48738 2546 48750
rect 9662 48802 9714 48814
rect 9662 48738 9714 48750
rect 13470 48802 13522 48814
rect 13470 48738 13522 48750
rect 14814 48802 14866 48814
rect 14814 48738 14866 48750
rect 16158 48802 16210 48814
rect 16158 48738 16210 48750
rect 18398 48802 18450 48814
rect 18398 48738 18450 48750
rect 18846 48802 18898 48814
rect 18846 48738 18898 48750
rect 20190 48802 20242 48814
rect 20190 48738 20242 48750
rect 22430 48802 22482 48814
rect 22430 48738 22482 48750
rect 23214 48802 23266 48814
rect 23214 48738 23266 48750
rect 32958 48802 33010 48814
rect 32958 48738 33010 48750
rect 33294 48802 33346 48814
rect 33294 48738 33346 48750
rect 33854 48802 33906 48814
rect 33854 48738 33906 48750
rect 34414 48802 34466 48814
rect 34414 48738 34466 48750
rect 34638 48802 34690 48814
rect 34638 48738 34690 48750
rect 36094 48802 36146 48814
rect 36094 48738 36146 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 3502 48466 3554 48478
rect 3502 48402 3554 48414
rect 16270 48466 16322 48478
rect 16270 48402 16322 48414
rect 16718 48466 16770 48478
rect 16718 48402 16770 48414
rect 17950 48466 18002 48478
rect 30494 48466 30546 48478
rect 19954 48414 19966 48466
rect 20018 48414 20030 48466
rect 17950 48402 18002 48414
rect 30494 48402 30546 48414
rect 31390 48466 31442 48478
rect 31390 48402 31442 48414
rect 38782 48466 38834 48478
rect 38782 48402 38834 48414
rect 7086 48354 7138 48366
rect 12126 48354 12178 48366
rect 10546 48302 10558 48354
rect 10610 48302 10622 48354
rect 7086 48290 7138 48302
rect 12126 48290 12178 48302
rect 15710 48354 15762 48366
rect 15710 48290 15762 48302
rect 17502 48354 17554 48366
rect 21534 48354 21586 48366
rect 19170 48302 19182 48354
rect 19234 48302 19246 48354
rect 19842 48302 19854 48354
rect 19906 48302 19918 48354
rect 17502 48290 17554 48302
rect 21534 48290 21586 48302
rect 21870 48354 21922 48366
rect 21870 48290 21922 48302
rect 22878 48354 22930 48366
rect 22878 48290 22930 48302
rect 23438 48354 23490 48366
rect 23438 48290 23490 48302
rect 23886 48354 23938 48366
rect 23886 48290 23938 48302
rect 23998 48354 24050 48366
rect 23998 48290 24050 48302
rect 26462 48354 26514 48366
rect 29822 48354 29874 48366
rect 31726 48354 31778 48366
rect 27346 48302 27358 48354
rect 27410 48302 27422 48354
rect 30818 48302 30830 48354
rect 30882 48302 30894 48354
rect 39106 48302 39118 48354
rect 39170 48302 39182 48354
rect 26462 48290 26514 48302
rect 29822 48290 29874 48302
rect 31726 48290 31778 48302
rect 6638 48242 6690 48254
rect 6638 48178 6690 48190
rect 7198 48242 7250 48254
rect 7198 48178 7250 48190
rect 9662 48242 9714 48254
rect 13582 48242 13634 48254
rect 10658 48190 10670 48242
rect 10722 48190 10734 48242
rect 11330 48190 11342 48242
rect 11394 48190 11406 48242
rect 11778 48190 11790 48242
rect 11842 48190 11854 48242
rect 9662 48178 9714 48190
rect 13582 48178 13634 48190
rect 13806 48242 13858 48254
rect 13806 48178 13858 48190
rect 14478 48242 14530 48254
rect 14478 48178 14530 48190
rect 15374 48242 15426 48254
rect 20078 48242 20130 48254
rect 18050 48190 18062 48242
rect 18114 48190 18126 48242
rect 15374 48178 15426 48190
rect 20078 48178 20130 48190
rect 22766 48242 22818 48254
rect 22766 48178 22818 48190
rect 23102 48242 23154 48254
rect 23102 48178 23154 48190
rect 23326 48242 23378 48254
rect 23326 48178 23378 48190
rect 23662 48242 23714 48254
rect 23662 48178 23714 48190
rect 24558 48242 24610 48254
rect 24558 48178 24610 48190
rect 26574 48242 26626 48254
rect 31166 48242 31218 48254
rect 27122 48190 27134 48242
rect 27186 48190 27198 48242
rect 28690 48190 28702 48242
rect 28754 48190 28766 48242
rect 29026 48190 29038 48242
rect 29090 48190 29102 48242
rect 26574 48178 26626 48190
rect 31166 48178 31218 48190
rect 31502 48242 31554 48254
rect 33618 48190 33630 48242
rect 33682 48190 33694 48242
rect 31502 48178 31554 48190
rect 4062 48130 4114 48142
rect 4062 48066 4114 48078
rect 6078 48130 6130 48142
rect 6078 48066 6130 48078
rect 10222 48130 10274 48142
rect 10222 48066 10274 48078
rect 13358 48130 13410 48142
rect 20526 48130 20578 48142
rect 15250 48078 15262 48130
rect 15314 48078 15326 48130
rect 18274 48078 18286 48130
rect 18338 48078 18350 48130
rect 13358 48066 13410 48078
rect 20526 48066 20578 48078
rect 22430 48130 22482 48142
rect 22430 48066 22482 48078
rect 32174 48130 32226 48142
rect 39678 48130 39730 48142
rect 38210 48078 38222 48130
rect 38274 48078 38286 48130
rect 32174 48066 32226 48078
rect 39678 48066 39730 48078
rect 7086 48018 7138 48030
rect 7086 47954 7138 47966
rect 14030 48018 14082 48030
rect 14030 47954 14082 47966
rect 17390 48018 17442 48030
rect 23998 48018 24050 48030
rect 22194 47966 22206 48018
rect 22258 48015 22270 48018
rect 22530 48015 22542 48018
rect 22258 47969 22542 48015
rect 22258 47966 22270 47969
rect 22530 47966 22542 47969
rect 22594 47966 22606 48018
rect 17390 47954 17442 47966
rect 23998 47954 24050 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 3278 47682 3330 47694
rect 3278 47618 3330 47630
rect 18622 47682 18674 47694
rect 18622 47618 18674 47630
rect 3054 47570 3106 47582
rect 3054 47506 3106 47518
rect 8766 47570 8818 47582
rect 8766 47506 8818 47518
rect 28254 47570 28306 47582
rect 28254 47506 28306 47518
rect 32062 47570 32114 47582
rect 32062 47506 32114 47518
rect 33070 47570 33122 47582
rect 33070 47506 33122 47518
rect 35646 47570 35698 47582
rect 40002 47518 40014 47570
rect 40066 47518 40078 47570
rect 35646 47506 35698 47518
rect 2158 47458 2210 47470
rect 2158 47394 2210 47406
rect 2718 47458 2770 47470
rect 2718 47394 2770 47406
rect 3950 47458 4002 47470
rect 7870 47458 7922 47470
rect 14926 47458 14978 47470
rect 6626 47406 6638 47458
rect 6690 47406 6702 47458
rect 8306 47406 8318 47458
rect 8370 47406 8382 47458
rect 10658 47406 10670 47458
rect 10722 47406 10734 47458
rect 11106 47406 11118 47458
rect 11170 47406 11182 47458
rect 3950 47394 4002 47406
rect 7870 47394 7922 47406
rect 14926 47394 14978 47406
rect 15262 47458 15314 47470
rect 15262 47394 15314 47406
rect 17166 47458 17218 47470
rect 17166 47394 17218 47406
rect 18286 47458 18338 47470
rect 18286 47394 18338 47406
rect 18398 47458 18450 47470
rect 18398 47394 18450 47406
rect 19182 47458 19234 47470
rect 33742 47458 33794 47470
rect 20066 47406 20078 47458
rect 20130 47406 20142 47458
rect 20290 47406 20302 47458
rect 20354 47406 20366 47458
rect 25554 47406 25566 47458
rect 25618 47406 25630 47458
rect 27458 47406 27470 47458
rect 27522 47406 27534 47458
rect 29586 47406 29598 47458
rect 29650 47406 29662 47458
rect 30930 47406 30942 47458
rect 30994 47406 31006 47458
rect 31266 47406 31278 47458
rect 31330 47406 31342 47458
rect 19182 47394 19234 47406
rect 33742 47394 33794 47406
rect 34862 47458 34914 47470
rect 34862 47394 34914 47406
rect 35198 47458 35250 47470
rect 35198 47394 35250 47406
rect 38110 47458 38162 47470
rect 39006 47458 39058 47470
rect 38546 47406 38558 47458
rect 38610 47406 38622 47458
rect 42802 47406 42814 47458
rect 42866 47406 42878 47458
rect 38110 47394 38162 47406
rect 39006 47394 39058 47406
rect 4510 47346 4562 47358
rect 4510 47282 4562 47294
rect 6190 47346 6242 47358
rect 6190 47282 6242 47294
rect 7310 47346 7362 47358
rect 14030 47346 14082 47358
rect 9202 47294 9214 47346
rect 9266 47294 9278 47346
rect 12786 47294 12798 47346
rect 12850 47294 12862 47346
rect 7310 47282 7362 47294
rect 14030 47282 14082 47294
rect 17278 47346 17330 47358
rect 17278 47282 17330 47294
rect 18734 47346 18786 47358
rect 18734 47282 18786 47294
rect 19406 47346 19458 47358
rect 19406 47282 19458 47294
rect 19854 47346 19906 47358
rect 34638 47346 34690 47358
rect 25778 47294 25790 47346
rect 25842 47294 25854 47346
rect 27794 47294 27806 47346
rect 27858 47294 27870 47346
rect 29138 47294 29150 47346
rect 29202 47294 29214 47346
rect 33394 47294 33406 47346
rect 33458 47294 33470 47346
rect 42130 47294 42142 47346
rect 42194 47294 42206 47346
rect 19854 47282 19906 47294
rect 34638 47282 34690 47294
rect 15038 47234 15090 47246
rect 3602 47182 3614 47234
rect 3666 47182 3678 47234
rect 10098 47182 10110 47234
rect 10162 47182 10174 47234
rect 15038 47170 15090 47182
rect 16494 47234 16546 47246
rect 16494 47170 16546 47182
rect 17502 47234 17554 47246
rect 17502 47170 17554 47182
rect 19294 47234 19346 47246
rect 19294 47170 19346 47182
rect 19742 47234 19794 47246
rect 19742 47170 19794 47182
rect 35086 47234 35138 47246
rect 39454 47234 39506 47246
rect 38770 47182 38782 47234
rect 38834 47182 38846 47234
rect 35086 47170 35138 47182
rect 39454 47170 39506 47182
rect 39566 47234 39618 47246
rect 39566 47170 39618 47182
rect 39678 47234 39730 47246
rect 39678 47170 39730 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 2494 46898 2546 46910
rect 2494 46834 2546 46846
rect 13694 46898 13746 46910
rect 13694 46834 13746 46846
rect 16158 46898 16210 46910
rect 16158 46834 16210 46846
rect 32622 46898 32674 46910
rect 32622 46834 32674 46846
rect 34078 46898 34130 46910
rect 34078 46834 34130 46846
rect 38446 46898 38498 46910
rect 38446 46834 38498 46846
rect 40350 46898 40402 46910
rect 40350 46834 40402 46846
rect 41358 46898 41410 46910
rect 41358 46834 41410 46846
rect 1710 46786 1762 46798
rect 1710 46722 1762 46734
rect 2046 46786 2098 46798
rect 2046 46722 2098 46734
rect 2942 46786 2994 46798
rect 6414 46786 6466 46798
rect 3714 46734 3726 46786
rect 3778 46734 3790 46786
rect 4834 46734 4846 46786
rect 4898 46734 4910 46786
rect 2942 46722 2994 46734
rect 6414 46722 6466 46734
rect 7870 46786 7922 46798
rect 13134 46786 13186 46798
rect 15710 46786 15762 46798
rect 33518 46786 33570 46798
rect 38782 46786 38834 46798
rect 40910 46786 40962 46798
rect 10322 46734 10334 46786
rect 10386 46734 10398 46786
rect 11330 46734 11342 46786
rect 11394 46734 11406 46786
rect 13346 46734 13358 46786
rect 13410 46734 13422 46786
rect 20738 46734 20750 46786
rect 20802 46734 20814 46786
rect 22642 46734 22654 46786
rect 22706 46734 22718 46786
rect 30146 46734 30158 46786
rect 30210 46734 30222 46786
rect 36642 46734 36654 46786
rect 36706 46734 36718 46786
rect 39442 46734 39454 46786
rect 39506 46734 39518 46786
rect 7870 46722 7922 46734
rect 13134 46722 13186 46734
rect 15710 46722 15762 46734
rect 33518 46722 33570 46734
rect 38782 46722 38834 46734
rect 40910 46722 40962 46734
rect 41134 46786 41186 46798
rect 41134 46722 41186 46734
rect 4510 46674 4562 46686
rect 7310 46674 7362 46686
rect 15038 46674 15090 46686
rect 23102 46674 23154 46686
rect 3938 46622 3950 46674
rect 4002 46622 4014 46674
rect 6962 46622 6974 46674
rect 7026 46622 7038 46674
rect 10770 46622 10782 46674
rect 10834 46622 10846 46674
rect 11442 46622 11454 46674
rect 11506 46622 11518 46674
rect 14690 46622 14702 46674
rect 14754 46622 14766 46674
rect 21298 46622 21310 46674
rect 21362 46622 21374 46674
rect 21522 46622 21534 46674
rect 21586 46622 21598 46674
rect 22082 46622 22094 46674
rect 22146 46622 22158 46674
rect 4510 46610 4562 46622
rect 7310 46610 7362 46622
rect 15038 46610 15090 46622
rect 23102 46610 23154 46622
rect 24222 46674 24274 46686
rect 33070 46674 33122 46686
rect 25218 46622 25230 46674
rect 25282 46622 25294 46674
rect 24222 46610 24274 46622
rect 33070 46610 33122 46622
rect 33294 46674 33346 46686
rect 33294 46610 33346 46622
rect 33742 46674 33794 46686
rect 39118 46674 39170 46686
rect 37314 46622 37326 46674
rect 37378 46622 37390 46674
rect 33742 46610 33794 46622
rect 39118 46610 39170 46622
rect 41470 46674 41522 46686
rect 41470 46610 41522 46622
rect 23662 46562 23714 46574
rect 3826 46510 3838 46562
rect 3890 46510 3902 46562
rect 5954 46510 5966 46562
rect 6018 46510 6030 46562
rect 14354 46510 14366 46562
rect 14418 46510 14430 46562
rect 22418 46510 22430 46562
rect 22482 46510 22494 46562
rect 23662 46498 23714 46510
rect 24782 46562 24834 46574
rect 34514 46510 34526 46562
rect 34578 46510 34590 46562
rect 24782 46498 24834 46510
rect 3054 46450 3106 46462
rect 38670 46450 38722 46462
rect 15026 46398 15038 46450
rect 15090 46398 15102 46450
rect 3054 46386 3106 46398
rect 38670 46386 38722 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 33630 46114 33682 46126
rect 33630 46050 33682 46062
rect 9886 46002 9938 46014
rect 9886 45938 9938 45950
rect 14478 46002 14530 46014
rect 14478 45938 14530 45950
rect 17726 46002 17778 46014
rect 17726 45938 17778 45950
rect 22206 46002 22258 46014
rect 32062 46002 32114 46014
rect 26898 45950 26910 46002
rect 26962 45950 26974 46002
rect 22206 45938 22258 45950
rect 32062 45938 32114 45950
rect 32846 46002 32898 46014
rect 34414 46002 34466 46014
rect 33954 45950 33966 46002
rect 34018 45950 34030 46002
rect 32846 45938 32898 45950
rect 34414 45938 34466 45950
rect 41022 46002 41074 46014
rect 41022 45938 41074 45950
rect 3950 45890 4002 45902
rect 7198 45890 7250 45902
rect 8654 45890 8706 45902
rect 12126 45890 12178 45902
rect 6850 45838 6862 45890
rect 6914 45838 6926 45890
rect 7634 45838 7646 45890
rect 7698 45838 7710 45890
rect 10322 45838 10334 45890
rect 10386 45838 10398 45890
rect 3950 45826 4002 45838
rect 7198 45826 7250 45838
rect 8654 45826 8706 45838
rect 12126 45826 12178 45838
rect 13918 45890 13970 45902
rect 13918 45826 13970 45838
rect 15934 45890 15986 45902
rect 17278 45890 17330 45902
rect 16370 45838 16382 45890
rect 16434 45838 16446 45890
rect 16706 45838 16718 45890
rect 16770 45838 16782 45890
rect 15934 45826 15986 45838
rect 17278 45826 17330 45838
rect 19966 45890 20018 45902
rect 19966 45826 20018 45838
rect 20078 45890 20130 45902
rect 21982 45890 22034 45902
rect 21522 45838 21534 45890
rect 21586 45838 21598 45890
rect 20078 45826 20130 45838
rect 21982 45826 22034 45838
rect 24446 45890 24498 45902
rect 32734 45890 32786 45902
rect 24770 45838 24782 45890
rect 24834 45838 24846 45890
rect 26786 45838 26798 45890
rect 26850 45838 26862 45890
rect 29362 45838 29374 45890
rect 29426 45838 29438 45890
rect 30930 45838 30942 45890
rect 30994 45838 31006 45890
rect 31826 45838 31838 45890
rect 31890 45838 31902 45890
rect 24446 45826 24498 45838
rect 32734 45826 32786 45838
rect 32958 45890 33010 45902
rect 32958 45826 33010 45838
rect 34526 45890 34578 45902
rect 34526 45826 34578 45838
rect 41582 45890 41634 45902
rect 41582 45826 41634 45838
rect 41918 45890 41970 45902
rect 41918 45826 41970 45838
rect 1710 45778 1762 45790
rect 1710 45714 1762 45726
rect 4510 45778 4562 45790
rect 4510 45714 4562 45726
rect 6526 45778 6578 45790
rect 6526 45714 6578 45726
rect 9326 45778 9378 45790
rect 9326 45714 9378 45726
rect 10894 45788 10946 45800
rect 10894 45724 10946 45736
rect 16158 45778 16210 45790
rect 22430 45778 22482 45790
rect 24558 45778 24610 45790
rect 27358 45778 27410 45790
rect 33182 45778 33234 45790
rect 21746 45726 21758 45778
rect 21810 45726 21822 45778
rect 23650 45726 23662 45778
rect 23714 45726 23726 45778
rect 24210 45726 24222 45778
rect 24274 45726 24286 45778
rect 24882 45726 24894 45778
rect 24946 45726 24958 45778
rect 29250 45726 29262 45778
rect 29314 45726 29326 45778
rect 16158 45714 16210 45726
rect 22430 45714 22482 45726
rect 24558 45714 24610 45726
rect 27358 45714 27410 45726
rect 33182 45714 33234 45726
rect 34750 45778 34802 45790
rect 34750 45714 34802 45726
rect 41358 45778 41410 45790
rect 41358 45714 41410 45726
rect 2046 45666 2098 45678
rect 2046 45602 2098 45614
rect 2494 45666 2546 45678
rect 2494 45602 2546 45614
rect 6638 45666 6690 45678
rect 6638 45602 6690 45614
rect 8094 45666 8146 45678
rect 8094 45602 8146 45614
rect 10446 45666 10498 45678
rect 10446 45602 10498 45614
rect 16046 45666 16098 45678
rect 16046 45602 16098 45614
rect 19742 45666 19794 45678
rect 19742 45602 19794 45614
rect 20638 45666 20690 45678
rect 20638 45602 20690 45614
rect 22542 45666 22594 45678
rect 22542 45602 22594 45614
rect 33854 45666 33906 45678
rect 33854 45602 33906 45614
rect 34302 45666 34354 45678
rect 34302 45602 34354 45614
rect 38670 45666 38722 45678
rect 38670 45602 38722 45614
rect 41806 45666 41858 45678
rect 41806 45602 41858 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 2606 45330 2658 45342
rect 2606 45266 2658 45278
rect 3166 45330 3218 45342
rect 3166 45266 3218 45278
rect 8206 45330 8258 45342
rect 8206 45266 8258 45278
rect 11230 45330 11282 45342
rect 21422 45330 21474 45342
rect 39230 45330 39282 45342
rect 19730 45278 19742 45330
rect 19794 45278 19806 45330
rect 21634 45278 21646 45330
rect 21698 45278 21710 45330
rect 23314 45278 23326 45330
rect 23378 45278 23390 45330
rect 27570 45278 27582 45330
rect 27634 45278 27646 45330
rect 11230 45266 11282 45278
rect 21422 45266 21474 45278
rect 39230 45266 39282 45278
rect 7982 45218 8034 45230
rect 7982 45154 8034 45166
rect 10670 45218 10722 45230
rect 22318 45218 22370 45230
rect 28702 45218 28754 45230
rect 19058 45166 19070 45218
rect 19122 45166 19134 45218
rect 19394 45166 19406 45218
rect 19458 45166 19470 45218
rect 26226 45166 26238 45218
rect 26290 45166 26302 45218
rect 10670 45154 10722 45166
rect 22318 45154 22370 45166
rect 28702 45154 28754 45166
rect 39006 45218 39058 45230
rect 39006 45154 39058 45166
rect 39342 45218 39394 45230
rect 42354 45166 42366 45218
rect 42418 45166 42430 45218
rect 39342 45154 39394 45166
rect 2494 45106 2546 45118
rect 2494 45042 2546 45054
rect 3054 45106 3106 45118
rect 6862 45106 6914 45118
rect 7758 45106 7810 45118
rect 4162 45054 4174 45106
rect 4226 45054 4238 45106
rect 6962 45054 6974 45106
rect 7026 45054 7038 45106
rect 3054 45042 3106 45054
rect 6862 45042 6914 45054
rect 7758 45042 7810 45054
rect 9774 45106 9826 45118
rect 9774 45042 9826 45054
rect 13694 45106 13746 45118
rect 13694 45042 13746 45054
rect 19966 45106 20018 45118
rect 19966 45042 20018 45054
rect 20750 45106 20802 45118
rect 20750 45042 20802 45054
rect 22094 45106 22146 45118
rect 22094 45042 22146 45054
rect 22206 45106 22258 45118
rect 22206 45042 22258 45054
rect 22766 45106 22818 45118
rect 29822 45106 29874 45118
rect 26114 45054 26126 45106
rect 26178 45054 26190 45106
rect 22766 45042 22818 45054
rect 29822 45042 29874 45054
rect 32510 45106 32562 45118
rect 39566 45106 39618 45118
rect 33394 45054 33406 45106
rect 33458 45054 33470 45106
rect 41570 45054 41582 45106
rect 41634 45054 41646 45106
rect 32510 45042 32562 45054
rect 39566 45042 39618 45054
rect 3726 44994 3778 45006
rect 11454 44994 11506 45006
rect 6738 44942 6750 44994
rect 6802 44942 6814 44994
rect 8194 44942 8206 44994
rect 8258 44942 8270 44994
rect 3726 44930 3778 44942
rect 11454 44930 11506 44942
rect 14254 44994 14306 45006
rect 14254 44930 14306 44942
rect 18622 44994 18674 45006
rect 18622 44930 18674 44942
rect 20302 44994 20354 45006
rect 20302 44930 20354 44942
rect 20526 44994 20578 45006
rect 20526 44930 20578 44942
rect 24670 44994 24722 45006
rect 24670 44930 24722 44942
rect 25342 44994 25394 45006
rect 25342 44930 25394 44942
rect 25790 44994 25842 45006
rect 25790 44930 25842 44942
rect 30382 44994 30434 45006
rect 37090 44942 37102 44994
rect 37154 44942 37166 44994
rect 44482 44942 44494 44994
rect 44546 44942 44558 44994
rect 30382 44930 30434 44942
rect 2606 44882 2658 44894
rect 2606 44818 2658 44830
rect 3166 44882 3218 44894
rect 3166 44818 3218 44830
rect 20974 44882 21026 44894
rect 20974 44818 21026 44830
rect 22990 44882 23042 44894
rect 22990 44818 23042 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 17278 44546 17330 44558
rect 17278 44482 17330 44494
rect 26014 44546 26066 44558
rect 26014 44482 26066 44494
rect 29934 44546 29986 44558
rect 29934 44482 29986 44494
rect 34526 44546 34578 44558
rect 34526 44482 34578 44494
rect 12574 44434 12626 44446
rect 8530 44382 8542 44434
rect 8594 44382 8606 44434
rect 10098 44382 10110 44434
rect 10162 44382 10174 44434
rect 12574 44370 12626 44382
rect 14814 44434 14866 44446
rect 14814 44370 14866 44382
rect 16158 44434 16210 44446
rect 33518 44434 33570 44446
rect 17602 44382 17614 44434
rect 17666 44382 17678 44434
rect 23426 44382 23438 44434
rect 23490 44382 23502 44434
rect 25778 44382 25790 44434
rect 25842 44382 25854 44434
rect 27794 44382 27806 44434
rect 27858 44382 27870 44434
rect 16158 44370 16210 44382
rect 33518 44370 33570 44382
rect 35422 44434 35474 44446
rect 41134 44434 41186 44446
rect 37202 44382 37214 44434
rect 37266 44382 37278 44434
rect 39330 44382 39342 44434
rect 39394 44382 39406 44434
rect 35422 44370 35474 44382
rect 41134 44370 41186 44382
rect 10222 44322 10274 44334
rect 11342 44322 11394 44334
rect 15710 44322 15762 44334
rect 6850 44270 6862 44322
rect 6914 44270 6926 44322
rect 10994 44270 11006 44322
rect 11058 44270 11070 44322
rect 11554 44270 11566 44322
rect 11618 44270 11630 44322
rect 12786 44270 12798 44322
rect 12850 44270 12862 44322
rect 14354 44270 14366 44322
rect 14418 44270 14430 44322
rect 15250 44270 15262 44322
rect 15314 44270 15326 44322
rect 10222 44258 10274 44270
rect 11342 44258 11394 44270
rect 15710 44258 15762 44270
rect 16382 44322 16434 44334
rect 16382 44258 16434 44270
rect 16606 44322 16658 44334
rect 16606 44258 16658 44270
rect 16830 44322 16882 44334
rect 26238 44322 26290 44334
rect 18386 44270 18398 44322
rect 18450 44270 18462 44322
rect 19058 44270 19070 44322
rect 19122 44270 19134 44322
rect 23090 44270 23102 44322
rect 23154 44270 23166 44322
rect 25218 44270 25230 44322
rect 25282 44270 25294 44322
rect 16830 44258 16882 44270
rect 26238 44258 26290 44270
rect 26910 44322 26962 44334
rect 29150 44322 29202 44334
rect 40574 44322 40626 44334
rect 28130 44270 28142 44322
rect 28194 44270 28206 44322
rect 30818 44270 30830 44322
rect 30882 44270 30894 44322
rect 32386 44270 32398 44322
rect 32450 44270 32462 44322
rect 33282 44270 33294 44322
rect 33346 44270 33358 44322
rect 34178 44270 34190 44322
rect 34242 44270 34254 44322
rect 34738 44270 34750 44322
rect 34802 44270 34814 44322
rect 40002 44270 40014 44322
rect 40066 44270 40078 44322
rect 26910 44258 26962 44270
rect 29150 44258 29202 44270
rect 40574 44258 40626 44270
rect 41022 44322 41074 44334
rect 41022 44258 41074 44270
rect 8094 44210 8146 44222
rect 5730 44158 5742 44210
rect 5794 44158 5806 44210
rect 8094 44146 8146 44158
rect 10558 44210 10610 44222
rect 10558 44146 10610 44158
rect 12462 44210 12514 44222
rect 24782 44210 24834 44222
rect 26798 44210 26850 44222
rect 34974 44210 35026 44222
rect 18050 44158 18062 44210
rect 18114 44158 18126 44210
rect 19282 44158 19294 44210
rect 19346 44158 19358 44210
rect 25106 44158 25118 44210
rect 25170 44158 25182 44210
rect 26562 44158 26574 44210
rect 26626 44158 26638 44210
rect 30594 44158 30606 44210
rect 30658 44158 30670 44210
rect 12462 44146 12514 44158
rect 24782 44146 24834 44158
rect 26798 44146 26850 44158
rect 34974 44146 35026 44158
rect 13694 44098 13746 44110
rect 11778 44046 11790 44098
rect 11842 44046 11854 44098
rect 13694 44034 13746 44046
rect 21422 44098 21474 44110
rect 21422 44034 21474 44046
rect 22654 44098 22706 44110
rect 22654 44034 22706 44046
rect 24334 44098 24386 44110
rect 41246 44098 41298 44110
rect 34626 44046 34638 44098
rect 34690 44046 34702 44098
rect 24334 44034 24386 44046
rect 41246 44034 41298 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 17502 43762 17554 43774
rect 29598 43762 29650 43774
rect 22194 43710 22206 43762
rect 22258 43710 22270 43762
rect 17502 43698 17554 43710
rect 29598 43698 29650 43710
rect 39566 43762 39618 43774
rect 39566 43698 39618 43710
rect 41134 43762 41186 43774
rect 41134 43698 41186 43710
rect 3502 43650 3554 43662
rect 3502 43586 3554 43598
rect 5294 43650 5346 43662
rect 5294 43586 5346 43598
rect 6190 43650 6242 43662
rect 6190 43586 6242 43598
rect 6414 43650 6466 43662
rect 6414 43586 6466 43598
rect 7422 43650 7474 43662
rect 7422 43586 7474 43598
rect 11118 43650 11170 43662
rect 11118 43586 11170 43598
rect 17390 43650 17442 43662
rect 17390 43586 17442 43598
rect 17614 43650 17666 43662
rect 17614 43586 17666 43598
rect 17726 43650 17778 43662
rect 21646 43650 21698 43662
rect 17826 43598 17838 43650
rect 17890 43598 17902 43650
rect 18610 43598 18622 43650
rect 18674 43598 18686 43650
rect 17726 43586 17778 43598
rect 21646 43586 21698 43598
rect 26350 43650 26402 43662
rect 26350 43586 26402 43598
rect 27134 43650 27186 43662
rect 27134 43586 27186 43598
rect 29150 43650 29202 43662
rect 29150 43586 29202 43598
rect 30942 43650 30994 43662
rect 30942 43586 30994 43598
rect 31726 43650 31778 43662
rect 37438 43650 37490 43662
rect 32050 43598 32062 43650
rect 32114 43598 32126 43650
rect 33394 43598 33406 43650
rect 33458 43598 33470 43650
rect 34626 43598 34638 43650
rect 34690 43598 34702 43650
rect 31726 43586 31778 43598
rect 37438 43586 37490 43598
rect 38782 43650 38834 43662
rect 38782 43586 38834 43598
rect 39230 43650 39282 43662
rect 39230 43586 39282 43598
rect 39454 43650 39506 43662
rect 39454 43586 39506 43598
rect 39678 43650 39730 43662
rect 39678 43586 39730 43598
rect 41582 43650 41634 43662
rect 41582 43586 41634 43598
rect 2382 43538 2434 43550
rect 2382 43474 2434 43486
rect 2494 43538 2546 43550
rect 2494 43474 2546 43486
rect 2718 43538 2770 43550
rect 8766 43538 8818 43550
rect 2930 43486 2942 43538
rect 2994 43486 3006 43538
rect 4834 43486 4846 43538
rect 4898 43486 4910 43538
rect 6962 43486 6974 43538
rect 7026 43486 7038 43538
rect 8306 43486 8318 43538
rect 8370 43486 8382 43538
rect 2718 43474 2770 43486
rect 8766 43474 8818 43486
rect 9102 43538 9154 43550
rect 9102 43474 9154 43486
rect 9998 43538 10050 43550
rect 10894 43538 10946 43550
rect 10098 43486 10110 43538
rect 10162 43486 10174 43538
rect 9998 43474 10050 43486
rect 10894 43474 10946 43486
rect 12238 43538 12290 43550
rect 12238 43474 12290 43486
rect 13022 43538 13074 43550
rect 13022 43474 13074 43486
rect 13918 43538 13970 43550
rect 23438 43538 23490 43550
rect 18498 43486 18510 43538
rect 18562 43486 18574 43538
rect 20514 43486 20526 43538
rect 20578 43486 20590 43538
rect 13918 43474 13970 43486
rect 23438 43474 23490 43486
rect 23998 43538 24050 43550
rect 23998 43474 24050 43486
rect 24670 43538 24722 43550
rect 24670 43474 24722 43486
rect 25566 43538 25618 43550
rect 25566 43474 25618 43486
rect 25678 43538 25730 43550
rect 37326 43538 37378 43550
rect 25890 43486 25902 43538
rect 25954 43486 25966 43538
rect 26562 43486 26574 43538
rect 26626 43486 26638 43538
rect 28578 43486 28590 43538
rect 28642 43486 28654 43538
rect 33170 43486 33182 43538
rect 33234 43486 33246 43538
rect 33954 43486 33966 43538
rect 34018 43486 34030 43538
rect 25678 43474 25730 43486
rect 37326 43474 37378 43486
rect 41358 43538 41410 43550
rect 41358 43474 41410 43486
rect 1822 43426 1874 43438
rect 4062 43426 4114 43438
rect 2818 43374 2830 43426
rect 2882 43374 2894 43426
rect 1822 43362 1874 43374
rect 4062 43362 4114 43374
rect 4398 43426 4450 43438
rect 4398 43362 4450 43374
rect 5854 43426 5906 43438
rect 5854 43362 5906 43374
rect 6302 43426 6354 43438
rect 12350 43426 12402 43438
rect 7858 43374 7870 43426
rect 7922 43374 7934 43426
rect 10210 43374 10222 43426
rect 10274 43374 10286 43426
rect 6302 43362 6354 43374
rect 12350 43362 12402 43374
rect 12574 43426 12626 43438
rect 12574 43362 12626 43374
rect 14478 43426 14530 43438
rect 14478 43362 14530 43374
rect 23102 43426 23154 43438
rect 23102 43362 23154 43374
rect 25342 43426 25394 43438
rect 25342 43362 25394 43374
rect 32510 43426 32562 43438
rect 41246 43426 41298 43438
rect 36754 43374 36766 43426
rect 36818 43374 36830 43426
rect 32510 43362 32562 43374
rect 41246 43362 41298 43374
rect 30718 43314 30770 43326
rect 30718 43250 30770 43262
rect 31054 43314 31106 43326
rect 31054 43250 31106 43262
rect 38670 43314 38722 43326
rect 38670 43250 38722 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 24670 42978 24722 42990
rect 24670 42914 24722 42926
rect 28366 42978 28418 42990
rect 28366 42914 28418 42926
rect 28254 42866 28306 42878
rect 33854 42866 33906 42878
rect 13906 42814 13918 42866
rect 13970 42814 13982 42866
rect 21746 42814 21758 42866
rect 21810 42814 21822 42866
rect 25442 42814 25454 42866
rect 25506 42814 25518 42866
rect 30370 42814 30382 42866
rect 30434 42814 30446 42866
rect 28254 42802 28306 42814
rect 33854 42802 33906 42814
rect 34750 42866 34802 42878
rect 34750 42802 34802 42814
rect 7086 42754 7138 42766
rect 1810 42702 1822 42754
rect 1874 42702 1886 42754
rect 7086 42690 7138 42702
rect 7646 42754 7698 42766
rect 13470 42754 13522 42766
rect 8754 42702 8766 42754
rect 8818 42702 8830 42754
rect 10770 42702 10782 42754
rect 10834 42702 10846 42754
rect 7646 42690 7698 42702
rect 13470 42690 13522 42702
rect 17614 42754 17666 42766
rect 22542 42754 22594 42766
rect 29822 42754 29874 42766
rect 30718 42754 30770 42766
rect 40126 42754 40178 42766
rect 18050 42702 18062 42754
rect 18114 42702 18126 42754
rect 25666 42702 25678 42754
rect 25730 42702 25742 42754
rect 27010 42702 27022 42754
rect 27074 42702 27086 42754
rect 29922 42702 29934 42754
rect 29986 42702 29998 42754
rect 31154 42702 31166 42754
rect 31218 42702 31230 42754
rect 33506 42702 33518 42754
rect 33570 42702 33582 42754
rect 17614 42690 17666 42702
rect 22542 42690 22594 42702
rect 29822 42690 29874 42702
rect 30718 42690 30770 42702
rect 40126 42690 40178 42702
rect 40350 42754 40402 42766
rect 40350 42690 40402 42702
rect 40686 42754 40738 42766
rect 40686 42690 40738 42702
rect 41022 42754 41074 42766
rect 41022 42690 41074 42702
rect 2046 42642 2098 42654
rect 2046 42578 2098 42590
rect 2718 42642 2770 42654
rect 2718 42578 2770 42590
rect 2830 42642 2882 42654
rect 2830 42578 2882 42590
rect 9886 42642 9938 42654
rect 9886 42578 9938 42590
rect 11342 42642 11394 42654
rect 11342 42578 11394 42590
rect 24558 42642 24610 42654
rect 26226 42590 26238 42642
rect 26290 42590 26302 42642
rect 30930 42590 30942 42642
rect 30994 42590 31006 42642
rect 32946 42590 32958 42642
rect 33010 42590 33022 42642
rect 24558 42578 24610 42590
rect 3054 42530 3106 42542
rect 21310 42530 21362 42542
rect 10882 42478 10894 42530
rect 10946 42478 10958 42530
rect 3054 42466 3106 42478
rect 21310 42466 21362 42478
rect 23102 42530 23154 42542
rect 23102 42466 23154 42478
rect 23886 42530 23938 42542
rect 23886 42466 23938 42478
rect 24334 42530 24386 42542
rect 24334 42466 24386 42478
rect 24670 42530 24722 42542
rect 24670 42466 24722 42478
rect 40686 42530 40738 42542
rect 40686 42466 40738 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 3502 42194 3554 42206
rect 16718 42194 16770 42206
rect 29262 42194 29314 42206
rect 8866 42142 8878 42194
rect 8930 42142 8942 42194
rect 20962 42142 20974 42194
rect 21026 42142 21038 42194
rect 3502 42130 3554 42142
rect 16718 42130 16770 42142
rect 29262 42130 29314 42142
rect 33182 42194 33234 42206
rect 35522 42142 35534 42194
rect 35586 42142 35598 42194
rect 33182 42130 33234 42142
rect 2270 42082 2322 42094
rect 2270 42018 2322 42030
rect 6414 42082 6466 42094
rect 6414 42018 6466 42030
rect 8430 42082 8482 42094
rect 16606 42082 16658 42094
rect 11218 42030 11230 42082
rect 11282 42030 11294 42082
rect 12114 42030 12126 42082
rect 12178 42030 12190 42082
rect 8430 42018 8482 42030
rect 16606 42018 16658 42030
rect 17838 42082 17890 42094
rect 17838 42018 17890 42030
rect 17950 42082 18002 42094
rect 17950 42018 18002 42030
rect 20750 42082 20802 42094
rect 20750 42018 20802 42030
rect 26350 42082 26402 42094
rect 26350 42018 26402 42030
rect 28590 42082 28642 42094
rect 28590 42018 28642 42030
rect 30606 42082 30658 42094
rect 30606 42018 30658 42030
rect 34526 42082 34578 42094
rect 34526 42018 34578 42030
rect 35086 42082 35138 42094
rect 35086 42018 35138 42030
rect 1822 41970 1874 41982
rect 1822 41906 1874 41918
rect 2494 41970 2546 41982
rect 2494 41906 2546 41918
rect 2718 41970 2770 41982
rect 5294 41970 5346 41982
rect 2930 41918 2942 41970
rect 2994 41918 3006 41970
rect 2718 41906 2770 41918
rect 5294 41906 5346 41918
rect 7310 41970 7362 41982
rect 18622 41970 18674 41982
rect 10546 41918 10558 41970
rect 10610 41918 10622 41970
rect 12226 41918 12238 41970
rect 12290 41918 12302 41970
rect 18386 41918 18398 41970
rect 18450 41918 18462 41970
rect 7310 41906 7362 41918
rect 18622 41906 18674 41918
rect 19966 41970 20018 41982
rect 19966 41906 20018 41918
rect 20302 41970 20354 41982
rect 20302 41906 20354 41918
rect 20526 41970 20578 41982
rect 20526 41906 20578 41918
rect 20974 41970 21026 41982
rect 20974 41906 21026 41918
rect 21982 41970 22034 41982
rect 21982 41906 22034 41918
rect 22094 41970 22146 41982
rect 22094 41906 22146 41918
rect 22206 41970 22258 41982
rect 24782 41970 24834 41982
rect 22418 41918 22430 41970
rect 22482 41918 22494 41970
rect 22206 41906 22258 41918
rect 24782 41906 24834 41918
rect 25678 41970 25730 41982
rect 25678 41906 25730 41918
rect 26238 41970 26290 41982
rect 26238 41906 26290 41918
rect 26574 41970 26626 41982
rect 33966 41970 34018 41982
rect 29698 41918 29710 41970
rect 29762 41918 29774 41970
rect 30146 41918 30158 41970
rect 30210 41918 30222 41970
rect 35298 41918 35310 41970
rect 35362 41918 35374 41970
rect 35858 41918 35870 41970
rect 35922 41918 35934 41970
rect 40898 41918 40910 41970
rect 40962 41918 40974 41970
rect 26574 41906 26626 41918
rect 33966 41906 34018 41918
rect 2606 41858 2658 41870
rect 2606 41794 2658 41806
rect 4062 41858 4114 41870
rect 18846 41858 18898 41870
rect 13346 41806 13358 41858
rect 13410 41806 13422 41858
rect 4062 41794 4114 41806
rect 18846 41794 18898 41806
rect 21534 41858 21586 41870
rect 21534 41794 21586 41806
rect 22878 41858 22930 41870
rect 22878 41794 22930 41806
rect 23214 41858 23266 41870
rect 25902 41858 25954 41870
rect 25330 41806 25342 41858
rect 25394 41806 25406 41858
rect 23214 41794 23266 41806
rect 25902 41794 25954 41806
rect 26910 41858 26962 41870
rect 26910 41794 26962 41806
rect 27582 41858 27634 41870
rect 27582 41794 27634 41806
rect 32174 41858 32226 41870
rect 32174 41794 32226 41806
rect 36318 41858 36370 41870
rect 36318 41794 36370 41806
rect 40126 41858 40178 41870
rect 41682 41806 41694 41858
rect 41746 41806 41758 41858
rect 43810 41806 43822 41858
rect 43874 41806 43886 41858
rect 40126 41794 40178 41806
rect 16718 41746 16770 41758
rect 16718 41682 16770 41694
rect 17950 41746 18002 41758
rect 17950 41682 18002 41694
rect 18958 41746 19010 41758
rect 18958 41682 19010 41694
rect 34302 41746 34354 41758
rect 34302 41682 34354 41694
rect 34638 41746 34690 41758
rect 34638 41682 34690 41694
rect 35534 41746 35586 41758
rect 35534 41682 35586 41694
rect 40014 41746 40066 41758
rect 40014 41682 40066 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 12014 41410 12066 41422
rect 12014 41346 12066 41358
rect 13918 41410 13970 41422
rect 13918 41346 13970 41358
rect 14366 41410 14418 41422
rect 14366 41346 14418 41358
rect 21758 41410 21810 41422
rect 21758 41346 21810 41358
rect 21982 41410 22034 41422
rect 21982 41346 22034 41358
rect 22094 41410 22146 41422
rect 27122 41358 27134 41410
rect 27186 41407 27198 41410
rect 28018 41407 28030 41410
rect 27186 41361 28030 41407
rect 27186 41358 27198 41361
rect 28018 41358 28030 41361
rect 28082 41358 28094 41410
rect 30370 41358 30382 41410
rect 30434 41358 30446 41410
rect 35410 41358 35422 41410
rect 35474 41358 35486 41410
rect 22094 41346 22146 41358
rect 7646 41298 7698 41310
rect 22878 41298 22930 41310
rect 27806 41298 27858 41310
rect 9538 41246 9550 41298
rect 9602 41246 9614 41298
rect 18162 41246 18174 41298
rect 18226 41246 18238 41298
rect 24994 41246 25006 41298
rect 25058 41246 25070 41298
rect 7646 41234 7698 41246
rect 22878 41234 22930 41246
rect 27806 41234 27858 41246
rect 28142 41298 28194 41310
rect 28142 41234 28194 41246
rect 28590 41298 28642 41310
rect 36094 41298 36146 41310
rect 30146 41246 30158 41298
rect 30210 41246 30222 41298
rect 37762 41246 37774 41298
rect 37826 41246 37838 41298
rect 39890 41246 39902 41298
rect 39954 41246 39966 41298
rect 28590 41234 28642 41246
rect 36094 41234 36146 41246
rect 1710 41186 1762 41198
rect 9214 41186 9266 41198
rect 14142 41186 14194 41198
rect 19630 41186 19682 41198
rect 5842 41134 5854 41186
rect 5906 41134 5918 41186
rect 9314 41134 9326 41186
rect 9378 41134 9390 41186
rect 11890 41134 11902 41186
rect 11954 41134 11966 41186
rect 17154 41134 17166 41186
rect 17218 41134 17230 41186
rect 17602 41134 17614 41186
rect 17666 41134 17678 41186
rect 1710 41122 1762 41134
rect 9214 41122 9266 41134
rect 14142 41122 14194 41134
rect 19630 41122 19682 41134
rect 19966 41186 20018 41198
rect 19966 41122 20018 41134
rect 20862 41186 20914 41198
rect 20862 41122 20914 41134
rect 21422 41186 21474 41198
rect 21422 41122 21474 41134
rect 21534 41186 21586 41198
rect 29150 41186 29202 41198
rect 34862 41186 34914 41198
rect 23202 41134 23214 41186
rect 23266 41134 23278 41186
rect 24882 41134 24894 41186
rect 24946 41134 24958 41186
rect 29362 41134 29374 41186
rect 29426 41134 29438 41186
rect 30482 41134 30494 41186
rect 30546 41134 30558 41186
rect 31378 41134 31390 41186
rect 31442 41134 31454 41186
rect 32946 41134 32958 41186
rect 33010 41134 33022 41186
rect 33842 41134 33854 41186
rect 33906 41134 33918 41186
rect 21534 41122 21586 41134
rect 29150 41122 29202 41134
rect 34862 41122 34914 41134
rect 35198 41186 35250 41198
rect 35410 41134 35422 41186
rect 35474 41134 35486 41186
rect 36978 41134 36990 41186
rect 37042 41134 37054 41186
rect 35198 41122 35250 41134
rect 2046 41074 2098 41086
rect 2046 41010 2098 41022
rect 2382 41074 2434 41086
rect 2382 41010 2434 41022
rect 2718 41074 2770 41086
rect 2718 41010 2770 41022
rect 6862 41074 6914 41086
rect 13694 41074 13746 41086
rect 20526 41074 20578 41086
rect 35982 41074 36034 41086
rect 12114 41022 12126 41074
rect 12178 41022 12190 41074
rect 15698 41022 15710 41074
rect 15762 41022 15774 41074
rect 19394 41022 19406 41074
rect 19458 41022 19470 41074
rect 23762 41022 23774 41074
rect 23826 41022 23838 41074
rect 24770 41022 24782 41074
rect 24834 41022 24846 41074
rect 31154 41022 31166 41074
rect 31218 41022 31230 41074
rect 6862 41010 6914 41022
rect 13694 41010 13746 41022
rect 20526 41010 20578 41022
rect 35982 41010 36034 41022
rect 7310 40962 7362 40974
rect 14814 40962 14866 40974
rect 9650 40910 9662 40962
rect 9714 40910 9726 40962
rect 7310 40898 7362 40910
rect 14814 40898 14866 40910
rect 15150 40962 15202 40974
rect 15150 40898 15202 40910
rect 19854 40962 19906 40974
rect 19854 40898 19906 40910
rect 20638 40962 20690 40974
rect 20638 40898 20690 40910
rect 27246 40962 27298 40974
rect 35646 40962 35698 40974
rect 32946 40910 32958 40962
rect 33010 40910 33022 40962
rect 27246 40898 27298 40910
rect 35646 40898 35698 40910
rect 36206 40962 36258 40974
rect 36206 40898 36258 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 12350 40626 12402 40638
rect 12350 40562 12402 40574
rect 13134 40626 13186 40638
rect 18174 40626 18226 40638
rect 16370 40574 16382 40626
rect 16434 40574 16446 40626
rect 13134 40562 13186 40574
rect 18174 40562 18226 40574
rect 19518 40626 19570 40638
rect 19518 40562 19570 40574
rect 21086 40626 21138 40638
rect 21086 40562 21138 40574
rect 22654 40626 22706 40638
rect 22654 40562 22706 40574
rect 24110 40626 24162 40638
rect 24110 40562 24162 40574
rect 25678 40626 25730 40638
rect 27134 40626 27186 40638
rect 26674 40574 26686 40626
rect 26738 40574 26750 40626
rect 25678 40562 25730 40574
rect 27134 40562 27186 40574
rect 34078 40626 34130 40638
rect 34078 40562 34130 40574
rect 34526 40626 34578 40638
rect 34526 40562 34578 40574
rect 35758 40626 35810 40638
rect 35758 40562 35810 40574
rect 36318 40626 36370 40638
rect 36318 40562 36370 40574
rect 2046 40514 2098 40526
rect 2046 40450 2098 40462
rect 4734 40514 4786 40526
rect 4734 40450 4786 40462
rect 6190 40514 6242 40526
rect 11790 40514 11842 40526
rect 34974 40514 35026 40526
rect 9762 40462 9774 40514
rect 9826 40462 9838 40514
rect 15810 40462 15822 40514
rect 15874 40462 15886 40514
rect 16146 40462 16158 40514
rect 16210 40462 16222 40514
rect 17714 40462 17726 40514
rect 17778 40462 17790 40514
rect 18610 40462 18622 40514
rect 18674 40462 18686 40514
rect 6190 40450 6242 40462
rect 11790 40450 11842 40462
rect 34974 40450 35026 40462
rect 1710 40402 1762 40414
rect 1710 40338 1762 40350
rect 2494 40402 2546 40414
rect 2494 40338 2546 40350
rect 3390 40402 3442 40414
rect 3390 40338 3442 40350
rect 5294 40402 5346 40414
rect 5294 40338 5346 40350
rect 5742 40402 5794 40414
rect 9102 40402 9154 40414
rect 12910 40402 12962 40414
rect 8418 40350 8430 40402
rect 8482 40350 8494 40402
rect 8642 40350 8654 40402
rect 8706 40350 8718 40402
rect 9986 40350 9998 40402
rect 10050 40350 10062 40402
rect 5742 40338 5794 40350
rect 9102 40338 9154 40350
rect 12910 40338 12962 40350
rect 13582 40402 13634 40414
rect 14814 40402 14866 40414
rect 14354 40350 14366 40402
rect 14418 40350 14430 40402
rect 13582 40338 13634 40350
rect 14814 40338 14866 40350
rect 15374 40402 15426 40414
rect 15374 40338 15426 40350
rect 16606 40402 16658 40414
rect 18846 40402 18898 40414
rect 17490 40350 17502 40402
rect 17554 40350 17566 40402
rect 16606 40338 16658 40350
rect 18846 40338 18898 40350
rect 19294 40402 19346 40414
rect 19294 40338 19346 40350
rect 23102 40402 23154 40414
rect 23102 40338 23154 40350
rect 26126 40402 26178 40414
rect 35310 40402 35362 40414
rect 28242 40350 28254 40402
rect 28306 40350 28318 40402
rect 28802 40350 28814 40402
rect 28866 40350 28878 40402
rect 30482 40350 30494 40402
rect 30546 40350 30558 40402
rect 30818 40350 30830 40402
rect 30882 40350 30894 40402
rect 31154 40350 31166 40402
rect 31218 40350 31230 40402
rect 26126 40338 26178 40350
rect 35310 40338 35362 40350
rect 35422 40402 35474 40414
rect 35522 40350 35534 40402
rect 35586 40350 35598 40402
rect 35422 40338 35474 40350
rect 5406 40290 5458 40302
rect 12014 40290 12066 40302
rect 8754 40238 8766 40290
rect 8818 40238 8830 40290
rect 11330 40238 11342 40290
rect 11394 40238 11406 40290
rect 5406 40226 5458 40238
rect 12014 40226 12066 40238
rect 13022 40290 13074 40302
rect 13022 40226 13074 40238
rect 18510 40290 18562 40302
rect 18510 40226 18562 40238
rect 27806 40290 27858 40302
rect 36766 40290 36818 40302
rect 29810 40238 29822 40290
rect 29874 40238 29886 40290
rect 34626 40238 34638 40290
rect 34690 40238 34702 40290
rect 27806 40226 27858 40238
rect 36766 40226 36818 40238
rect 25342 40178 25394 40190
rect 23762 40126 23774 40178
rect 23826 40175 23838 40178
rect 24098 40175 24110 40178
rect 23826 40129 24110 40175
rect 23826 40126 23838 40129
rect 24098 40126 24110 40129
rect 24162 40126 24174 40178
rect 25342 40114 25394 40126
rect 25566 40178 25618 40190
rect 25566 40114 25618 40126
rect 25678 40178 25730 40190
rect 25678 40114 25730 40126
rect 26350 40178 26402 40190
rect 26350 40114 26402 40126
rect 34302 40178 34354 40190
rect 34302 40114 34354 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 7422 39842 7474 39854
rect 7422 39778 7474 39790
rect 28702 39842 28754 39854
rect 30258 39790 30270 39842
rect 30322 39790 30334 39842
rect 28702 39778 28754 39790
rect 6078 39730 6130 39742
rect 12686 39730 12738 39742
rect 11106 39678 11118 39730
rect 11170 39678 11182 39730
rect 6078 39666 6130 39678
rect 12686 39666 12738 39678
rect 22990 39730 23042 39742
rect 29598 39730 29650 39742
rect 26674 39678 26686 39730
rect 26738 39678 26750 39730
rect 32274 39678 32286 39730
rect 32338 39678 32350 39730
rect 22990 39666 23042 39678
rect 29598 39666 29650 39678
rect 3054 39618 3106 39630
rect 10670 39618 10722 39630
rect 14142 39618 14194 39630
rect 16382 39618 16434 39630
rect 27022 39618 27074 39630
rect 3938 39566 3950 39618
rect 4002 39566 4014 39618
rect 5058 39566 5070 39618
rect 5122 39566 5134 39618
rect 7970 39566 7982 39618
rect 8034 39566 8046 39618
rect 8642 39566 8654 39618
rect 8706 39566 8718 39618
rect 10770 39566 10782 39618
rect 10834 39566 10846 39618
rect 14914 39566 14926 39618
rect 14978 39566 14990 39618
rect 17378 39566 17390 39618
rect 17442 39566 17454 39618
rect 18722 39566 18734 39618
rect 18786 39566 18798 39618
rect 21298 39566 21310 39618
rect 21362 39566 21374 39618
rect 23314 39566 23326 39618
rect 23378 39566 23390 39618
rect 3054 39554 3106 39566
rect 10670 39554 10722 39566
rect 14142 39554 14194 39566
rect 16382 39554 16434 39566
rect 27022 39554 27074 39566
rect 27806 39618 27858 39630
rect 27806 39554 27858 39566
rect 28030 39618 28082 39630
rect 28030 39554 28082 39566
rect 28254 39618 28306 39630
rect 30718 39618 30770 39630
rect 30146 39566 30158 39618
rect 30210 39566 30222 39618
rect 28254 39554 28306 39566
rect 30718 39554 30770 39566
rect 30942 39618 30994 39630
rect 31378 39566 31390 39618
rect 31442 39566 31454 39618
rect 31826 39566 31838 39618
rect 31890 39566 31902 39618
rect 34066 39566 34078 39618
rect 34130 39566 34142 39618
rect 34962 39566 34974 39618
rect 35026 39566 35038 39618
rect 30942 39554 30994 39566
rect 2830 39506 2882 39518
rect 19630 39506 19682 39518
rect 23886 39506 23938 39518
rect 3378 39454 3390 39506
rect 3442 39454 3454 39506
rect 4946 39454 4958 39506
rect 5010 39454 5022 39506
rect 7858 39454 7870 39506
rect 7922 39454 7934 39506
rect 8754 39454 8766 39506
rect 8818 39454 8830 39506
rect 18162 39454 18174 39506
rect 18226 39454 18238 39506
rect 22418 39454 22430 39506
rect 22482 39454 22494 39506
rect 2830 39442 2882 39454
rect 19630 39442 19682 39454
rect 23886 39442 23938 39454
rect 25902 39506 25954 39518
rect 33842 39454 33854 39506
rect 33906 39454 33918 39506
rect 34738 39454 34750 39506
rect 34802 39454 34814 39506
rect 25902 39442 25954 39454
rect 2942 39394 2994 39406
rect 11566 39394 11618 39406
rect 3490 39342 3502 39394
rect 3554 39342 3566 39394
rect 2942 39330 2994 39342
rect 11566 39330 11618 39342
rect 14702 39394 14754 39406
rect 18050 39342 18062 39394
rect 18114 39342 18126 39394
rect 14702 39330 14754 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 3838 39058 3890 39070
rect 3838 38994 3890 39006
rect 4286 39058 4338 39070
rect 11790 39058 11842 39070
rect 15262 39058 15314 39070
rect 5730 39006 5742 39058
rect 5794 39006 5806 39058
rect 13010 39006 13022 39058
rect 13074 39006 13086 39058
rect 4286 38994 4338 39006
rect 11790 38994 11842 39006
rect 15262 38994 15314 39006
rect 19406 39058 19458 39070
rect 19406 38994 19458 39006
rect 21982 39058 22034 39070
rect 21982 38994 22034 39006
rect 22206 39058 22258 39070
rect 22206 38994 22258 39006
rect 23774 39058 23826 39070
rect 23774 38994 23826 39006
rect 24670 39058 24722 39070
rect 24670 38994 24722 39006
rect 25118 39058 25170 39070
rect 25118 38994 25170 39006
rect 27582 39058 27634 39070
rect 27582 38994 27634 39006
rect 29598 39058 29650 39070
rect 29598 38994 29650 39006
rect 15486 38946 15538 38958
rect 2370 38894 2382 38946
rect 2434 38894 2446 38946
rect 3490 38894 3502 38946
rect 3554 38894 3566 38946
rect 5618 38894 5630 38946
rect 5682 38894 5694 38946
rect 7074 38894 7086 38946
rect 7138 38894 7150 38946
rect 15486 38882 15538 38894
rect 24222 38946 24274 38958
rect 24222 38882 24274 38894
rect 26238 38946 26290 38958
rect 26238 38882 26290 38894
rect 26798 38946 26850 38958
rect 26798 38882 26850 38894
rect 28030 38946 28082 38958
rect 28030 38882 28082 38894
rect 30942 38946 30994 38958
rect 32386 38894 32398 38946
rect 32450 38894 32462 38946
rect 34290 38894 34302 38946
rect 34354 38894 34366 38946
rect 35522 38894 35534 38946
rect 35586 38894 35598 38946
rect 38210 38894 38222 38946
rect 38274 38894 38286 38946
rect 30942 38882 30994 38894
rect 5182 38834 5234 38846
rect 7646 38834 7698 38846
rect 2594 38782 2606 38834
rect 2658 38782 2670 38834
rect 6178 38782 6190 38834
rect 6242 38782 6254 38834
rect 6514 38782 6526 38834
rect 6578 38782 6590 38834
rect 5182 38770 5234 38782
rect 7646 38770 7698 38782
rect 7870 38834 7922 38846
rect 14478 38834 14530 38846
rect 12786 38782 12798 38834
rect 12850 38782 12862 38834
rect 14018 38782 14030 38834
rect 14082 38782 14094 38834
rect 7870 38770 7922 38782
rect 14478 38770 14530 38782
rect 14814 38834 14866 38846
rect 14814 38770 14866 38782
rect 15038 38834 15090 38846
rect 15038 38770 15090 38782
rect 20974 38834 21026 38846
rect 20974 38770 21026 38782
rect 21198 38834 21250 38846
rect 21198 38770 21250 38782
rect 21310 38834 21362 38846
rect 26014 38834 26066 38846
rect 21522 38782 21534 38834
rect 21586 38782 21598 38834
rect 21310 38770 21362 38782
rect 26014 38770 26066 38782
rect 26910 38834 26962 38846
rect 28366 38834 28418 38846
rect 36878 38834 36930 38846
rect 27122 38782 27134 38834
rect 27186 38782 27198 38834
rect 31266 38782 31278 38834
rect 31330 38782 31342 38834
rect 31714 38782 31726 38834
rect 31778 38782 31790 38834
rect 32498 38782 32510 38834
rect 32562 38782 32574 38834
rect 34962 38782 34974 38834
rect 35026 38782 35038 38834
rect 37426 38782 37438 38834
rect 37490 38782 37502 38834
rect 26910 38770 26962 38782
rect 28366 38770 28418 38782
rect 36878 38770 36930 38782
rect 1822 38722 1874 38734
rect 1822 38658 1874 38670
rect 7982 38722 8034 38734
rect 7982 38658 8034 38670
rect 8542 38722 8594 38734
rect 8542 38658 8594 38670
rect 12350 38722 12402 38734
rect 12350 38658 12402 38670
rect 18062 38722 18114 38734
rect 18062 38658 18114 38670
rect 18846 38722 18898 38734
rect 18846 38658 18898 38670
rect 19966 38722 20018 38734
rect 19966 38658 20018 38670
rect 20302 38722 20354 38734
rect 20302 38658 20354 38670
rect 22766 38722 22818 38734
rect 22766 38658 22818 38670
rect 23214 38722 23266 38734
rect 23214 38658 23266 38670
rect 25566 38722 25618 38734
rect 25566 38658 25618 38670
rect 26574 38722 26626 38734
rect 26574 38658 26626 38670
rect 28142 38722 28194 38734
rect 28142 38658 28194 38670
rect 28478 38722 28530 38734
rect 28478 38658 28530 38670
rect 29038 38722 29090 38734
rect 33842 38670 33854 38722
rect 33906 38670 33918 38722
rect 40338 38670 40350 38722
rect 40402 38670 40414 38722
rect 29038 38658 29090 38670
rect 7534 38610 7586 38622
rect 7534 38546 7586 38558
rect 15374 38610 15426 38622
rect 15374 38546 15426 38558
rect 25790 38610 25842 38622
rect 25790 38546 25842 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 4958 38274 5010 38286
rect 4958 38210 5010 38222
rect 13582 38274 13634 38286
rect 13582 38210 13634 38222
rect 19070 38274 19122 38286
rect 19070 38210 19122 38222
rect 20638 38274 20690 38286
rect 20638 38210 20690 38222
rect 19630 38162 19682 38174
rect 28366 38162 28418 38174
rect 7410 38110 7422 38162
rect 7474 38110 7486 38162
rect 11106 38110 11118 38162
rect 11170 38110 11182 38162
rect 12226 38110 12238 38162
rect 12290 38110 12302 38162
rect 15138 38110 15150 38162
rect 15202 38110 15214 38162
rect 27010 38110 27022 38162
rect 27074 38110 27086 38162
rect 19630 38098 19682 38110
rect 28366 38098 28418 38110
rect 29262 38162 29314 38174
rect 29262 38098 29314 38110
rect 30046 38162 30098 38174
rect 30046 38098 30098 38110
rect 32958 38162 33010 38174
rect 34290 38110 34302 38162
rect 34354 38110 34366 38162
rect 37202 38110 37214 38162
rect 37266 38110 37278 38162
rect 32958 38098 33010 38110
rect 2494 38050 2546 38062
rect 2494 37986 2546 37998
rect 3054 38050 3106 38062
rect 3054 37986 3106 37998
rect 4062 38050 4114 38062
rect 4062 37986 4114 37998
rect 4174 38050 4226 38062
rect 4174 37986 4226 37998
rect 4734 38050 4786 38062
rect 4734 37986 4786 37998
rect 5630 38050 5682 38062
rect 9550 38050 9602 38062
rect 11454 38050 11506 38062
rect 6514 37998 6526 38050
rect 6578 37998 6590 38050
rect 7746 37998 7758 38050
rect 7810 37998 7822 38050
rect 9986 37998 9998 38050
rect 10050 37998 10062 38050
rect 5630 37986 5682 37998
rect 9550 37986 9602 37998
rect 11454 37986 11506 37998
rect 11790 38050 11842 38062
rect 11790 37986 11842 37998
rect 11902 38050 11954 38062
rect 12798 38050 12850 38062
rect 12338 37998 12350 38050
rect 12402 37998 12414 38050
rect 11902 37986 11954 37998
rect 12798 37986 12850 37998
rect 14030 38050 14082 38062
rect 17278 38050 17330 38062
rect 15026 37998 15038 38050
rect 15090 37998 15102 38050
rect 15586 37998 15598 38050
rect 15650 37998 15662 38050
rect 14030 37986 14082 37998
rect 17278 37986 17330 37998
rect 17950 38050 18002 38062
rect 17950 37986 18002 37998
rect 18398 38050 18450 38062
rect 18398 37986 18450 37998
rect 18510 38050 18562 38062
rect 18510 37986 18562 37998
rect 18734 38050 18786 38062
rect 18734 37986 18786 37998
rect 18958 38050 19010 38062
rect 18958 37986 19010 37998
rect 19966 38050 20018 38062
rect 19966 37986 20018 37998
rect 20414 38050 20466 38062
rect 28254 38050 28306 38062
rect 29822 38050 29874 38062
rect 24098 37998 24110 38050
rect 24162 37998 24174 38050
rect 26114 37998 26126 38050
rect 26178 37998 26190 38050
rect 28578 37998 28590 38050
rect 28642 37998 28654 38050
rect 20414 37986 20466 37998
rect 28254 37986 28306 37998
rect 29822 37986 29874 37998
rect 30494 38050 30546 38062
rect 30494 37986 30546 37998
rect 31838 38050 31890 38062
rect 37774 38050 37826 38062
rect 33394 37998 33406 38050
rect 33458 37998 33470 38050
rect 31838 37986 31890 37998
rect 37774 37986 37826 37998
rect 37998 38050 38050 38062
rect 37998 37986 38050 37998
rect 38222 38050 38274 38062
rect 38222 37986 38274 37998
rect 1710 37938 1762 37950
rect 1710 37874 1762 37886
rect 2606 37938 2658 37950
rect 2606 37874 2658 37886
rect 4286 37938 4338 37950
rect 10894 37938 10946 37950
rect 6962 37886 6974 37938
rect 7026 37886 7038 37938
rect 4286 37874 4338 37886
rect 10894 37874 10946 37886
rect 13470 37938 13522 37950
rect 16942 37938 16994 37950
rect 14466 37886 14478 37938
rect 14530 37886 14542 37938
rect 13470 37874 13522 37886
rect 16942 37874 16994 37886
rect 17838 37938 17890 37950
rect 22430 37938 22482 37950
rect 19730 37886 19742 37938
rect 19794 37886 19806 37938
rect 17838 37874 17890 37886
rect 22430 37874 22482 37886
rect 25230 37938 25282 37950
rect 25230 37874 25282 37886
rect 26686 37938 26738 37950
rect 26686 37874 26738 37886
rect 30606 37938 30658 37950
rect 30606 37874 30658 37886
rect 32062 37938 32114 37950
rect 32062 37874 32114 37886
rect 32174 37938 32226 37950
rect 32174 37874 32226 37886
rect 38446 37938 38498 37950
rect 38446 37874 38498 37886
rect 2046 37826 2098 37838
rect 2046 37762 2098 37774
rect 2830 37826 2882 37838
rect 2830 37762 2882 37774
rect 3614 37826 3666 37838
rect 3614 37762 3666 37774
rect 6190 37826 6242 37838
rect 9214 37826 9266 37838
rect 6850 37774 6862 37826
rect 6914 37774 6926 37826
rect 6190 37762 6242 37774
rect 9214 37762 9266 37774
rect 10670 37826 10722 37838
rect 10670 37762 10722 37774
rect 11118 37826 11170 37838
rect 11118 37762 11170 37774
rect 12126 37826 12178 37838
rect 12126 37762 12178 37774
rect 13694 37826 13746 37838
rect 13694 37762 13746 37774
rect 13918 37826 13970 37838
rect 16382 37826 16434 37838
rect 15810 37774 15822 37826
rect 15874 37774 15886 37826
rect 13918 37762 13970 37774
rect 16382 37762 16434 37774
rect 17390 37826 17442 37838
rect 17390 37762 17442 37774
rect 17614 37826 17666 37838
rect 17614 37762 17666 37774
rect 21422 37826 21474 37838
rect 21422 37762 21474 37774
rect 21870 37826 21922 37838
rect 21870 37762 21922 37774
rect 22990 37826 23042 37838
rect 22990 37762 23042 37774
rect 23438 37826 23490 37838
rect 23438 37762 23490 37774
rect 23774 37826 23826 37838
rect 23774 37762 23826 37774
rect 29710 37826 29762 37838
rect 29710 37762 29762 37774
rect 33854 37826 33906 37838
rect 33854 37762 33906 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 2606 37490 2658 37502
rect 2606 37426 2658 37438
rect 6302 37490 6354 37502
rect 10558 37490 10610 37502
rect 8194 37438 8206 37490
rect 8258 37438 8270 37490
rect 6302 37426 6354 37438
rect 10558 37426 10610 37438
rect 12574 37490 12626 37502
rect 12574 37426 12626 37438
rect 13022 37490 13074 37502
rect 13022 37426 13074 37438
rect 15822 37490 15874 37502
rect 26686 37490 26738 37502
rect 17938 37438 17950 37490
rect 18002 37438 18014 37490
rect 24658 37438 24670 37490
rect 24722 37438 24734 37490
rect 15822 37426 15874 37438
rect 26686 37426 26738 37438
rect 28030 37490 28082 37502
rect 28030 37426 28082 37438
rect 29038 37490 29090 37502
rect 29038 37426 29090 37438
rect 29486 37490 29538 37502
rect 29486 37426 29538 37438
rect 29710 37490 29762 37502
rect 29710 37426 29762 37438
rect 32062 37490 32114 37502
rect 39902 37490 39954 37502
rect 39554 37438 39566 37490
rect 39618 37438 39630 37490
rect 32062 37426 32114 37438
rect 39902 37426 39954 37438
rect 2046 37378 2098 37390
rect 2046 37314 2098 37326
rect 2494 37378 2546 37390
rect 2494 37314 2546 37326
rect 8766 37378 8818 37390
rect 8766 37314 8818 37326
rect 9774 37378 9826 37390
rect 16270 37378 16322 37390
rect 12114 37326 12126 37378
rect 12178 37326 12190 37378
rect 9774 37314 9826 37326
rect 16270 37314 16322 37326
rect 16494 37378 16546 37390
rect 16494 37314 16546 37326
rect 18286 37378 18338 37390
rect 18286 37314 18338 37326
rect 18398 37378 18450 37390
rect 18398 37314 18450 37326
rect 19182 37378 19234 37390
rect 19182 37314 19234 37326
rect 19406 37378 19458 37390
rect 28254 37378 28306 37390
rect 23874 37326 23886 37378
rect 23938 37326 23950 37378
rect 25778 37326 25790 37378
rect 25842 37326 25854 37378
rect 26114 37326 26126 37378
rect 26178 37326 26190 37378
rect 19406 37314 19458 37326
rect 28254 37314 28306 37326
rect 29598 37378 29650 37390
rect 29598 37314 29650 37326
rect 32286 37378 32338 37390
rect 40350 37378 40402 37390
rect 35970 37326 35982 37378
rect 36034 37326 36046 37378
rect 32286 37314 32338 37326
rect 40350 37314 40402 37326
rect 1710 37266 1762 37278
rect 8654 37266 8706 37278
rect 9886 37266 9938 37278
rect 15374 37266 15426 37278
rect 7746 37214 7758 37266
rect 7810 37214 7822 37266
rect 8978 37214 8990 37266
rect 9042 37214 9054 37266
rect 10098 37214 10110 37266
rect 10162 37214 10174 37266
rect 11890 37214 11902 37266
rect 11954 37214 11966 37266
rect 1710 37202 1762 37214
rect 8654 37202 8706 37214
rect 9886 37202 9938 37214
rect 15374 37202 15426 37214
rect 15934 37266 15986 37278
rect 15934 37202 15986 37214
rect 17614 37266 17666 37278
rect 17614 37202 17666 37214
rect 18622 37266 18674 37278
rect 18622 37202 18674 37214
rect 19070 37266 19122 37278
rect 27582 37266 27634 37278
rect 20850 37214 20862 37266
rect 20914 37214 20926 37266
rect 21074 37214 21086 37266
rect 21138 37214 21150 37266
rect 21522 37214 21534 37266
rect 21586 37214 21598 37266
rect 22754 37214 22766 37266
rect 22818 37214 22830 37266
rect 24434 37214 24446 37266
rect 24498 37214 24510 37266
rect 26450 37214 26462 37266
rect 26514 37214 26526 37266
rect 19070 37202 19122 37214
rect 27582 37202 27634 37214
rect 28366 37266 28418 37278
rect 28366 37202 28418 37214
rect 29822 37266 29874 37278
rect 34302 37266 34354 37278
rect 30034 37214 30046 37266
rect 30098 37214 30110 37266
rect 31042 37214 31054 37266
rect 31106 37214 31118 37266
rect 31266 37214 31278 37266
rect 31330 37214 31342 37266
rect 31490 37214 31502 37266
rect 31554 37214 31566 37266
rect 29822 37202 29874 37214
rect 34302 37202 34354 37214
rect 34862 37266 34914 37278
rect 35298 37214 35310 37266
rect 35362 37214 35374 37266
rect 34862 37202 34914 37214
rect 3166 37154 3218 37166
rect 9550 37154 9602 37166
rect 7410 37102 7422 37154
rect 7474 37102 7486 37154
rect 3166 37090 3218 37102
rect 9550 37090 9602 37102
rect 14926 37154 14978 37166
rect 14926 37090 14978 37102
rect 25454 37154 25506 37166
rect 25454 37090 25506 37102
rect 27806 37154 27858 37166
rect 38110 37154 38162 37166
rect 31938 37102 31950 37154
rect 32002 37102 32014 37154
rect 27806 37090 27858 37102
rect 38110 37090 38162 37102
rect 2606 37042 2658 37054
rect 2606 36978 2658 36990
rect 15150 37042 15202 37054
rect 15150 36978 15202 36990
rect 16158 37042 16210 37054
rect 16158 36978 16210 36990
rect 27134 37042 27186 37054
rect 27134 36978 27186 36990
rect 27358 37042 27410 37054
rect 40238 37042 40290 37054
rect 30482 36990 30494 37042
rect 30546 36990 30558 37042
rect 27358 36978 27410 36990
rect 40238 36978 40290 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 14142 36706 14194 36718
rect 7186 36654 7198 36706
rect 7250 36654 7262 36706
rect 14142 36642 14194 36654
rect 18174 36706 18226 36718
rect 18722 36654 18734 36706
rect 18786 36703 18798 36706
rect 20066 36703 20078 36706
rect 18786 36657 20078 36703
rect 18786 36654 18798 36657
rect 20066 36654 20078 36657
rect 20130 36654 20142 36706
rect 18174 36642 18226 36654
rect 8206 36594 8258 36606
rect 3602 36542 3614 36594
rect 3666 36542 3678 36594
rect 7074 36542 7086 36594
rect 7138 36542 7150 36594
rect 8206 36530 8258 36542
rect 12910 36594 12962 36606
rect 12910 36530 12962 36542
rect 17502 36594 17554 36606
rect 17502 36530 17554 36542
rect 18846 36594 18898 36606
rect 18846 36530 18898 36542
rect 27582 36594 27634 36606
rect 27582 36530 27634 36542
rect 31726 36594 31778 36606
rect 34638 36594 34690 36606
rect 33282 36542 33294 36594
rect 33346 36542 33358 36594
rect 31726 36530 31778 36542
rect 34638 36530 34690 36542
rect 36990 36594 37042 36606
rect 38882 36542 38894 36594
rect 38946 36542 38958 36594
rect 36990 36530 37042 36542
rect 8654 36482 8706 36494
rect 2482 36430 2494 36482
rect 2546 36430 2558 36482
rect 2706 36430 2718 36482
rect 2770 36430 2782 36482
rect 3266 36430 3278 36482
rect 3330 36430 3342 36482
rect 5730 36430 5742 36482
rect 5794 36430 5806 36482
rect 8654 36418 8706 36430
rect 14366 36482 14418 36494
rect 20414 36482 20466 36494
rect 18050 36430 18062 36482
rect 18114 36430 18126 36482
rect 14366 36418 14418 36430
rect 20414 36418 20466 36430
rect 20750 36482 20802 36494
rect 28702 36482 28754 36494
rect 22530 36430 22542 36482
rect 22594 36430 22606 36482
rect 24098 36430 24110 36482
rect 24162 36430 24174 36482
rect 25778 36430 25790 36482
rect 25842 36430 25854 36482
rect 26002 36430 26014 36482
rect 26066 36430 26078 36482
rect 20750 36418 20802 36430
rect 28702 36418 28754 36430
rect 29710 36482 29762 36494
rect 32846 36482 32898 36494
rect 32162 36430 32174 36482
rect 32226 36430 32238 36482
rect 29710 36418 29762 36430
rect 32846 36418 32898 36430
rect 36318 36482 36370 36494
rect 39554 36430 39566 36482
rect 39618 36430 39630 36482
rect 36318 36418 36370 36430
rect 6750 36370 6802 36382
rect 1922 36318 1934 36370
rect 1986 36318 1998 36370
rect 3826 36318 3838 36370
rect 3890 36318 3902 36370
rect 5954 36318 5966 36370
rect 6018 36318 6030 36370
rect 6750 36306 6802 36318
rect 10446 36370 10498 36382
rect 10446 36306 10498 36318
rect 13806 36370 13858 36382
rect 13806 36306 13858 36318
rect 18286 36370 18338 36382
rect 18286 36306 18338 36318
rect 20190 36370 20242 36382
rect 28366 36370 28418 36382
rect 22866 36318 22878 36370
rect 22930 36318 22942 36370
rect 23986 36318 23998 36370
rect 24050 36318 24062 36370
rect 20190 36306 20242 36318
rect 28366 36306 28418 36318
rect 35422 36370 35474 36382
rect 35422 36306 35474 36318
rect 4286 36258 4338 36270
rect 4286 36194 4338 36206
rect 4846 36258 4898 36270
rect 4846 36194 4898 36206
rect 8990 36258 9042 36270
rect 8990 36194 9042 36206
rect 14030 36258 14082 36270
rect 14030 36194 14082 36206
rect 17838 36258 17890 36270
rect 17838 36194 17890 36206
rect 19406 36258 19458 36270
rect 19406 36194 19458 36206
rect 19742 36258 19794 36270
rect 19742 36194 19794 36206
rect 20638 36258 20690 36270
rect 20638 36194 20690 36206
rect 21534 36258 21586 36270
rect 21534 36194 21586 36206
rect 21982 36258 22034 36270
rect 28030 36258 28082 36270
rect 23874 36206 23886 36258
rect 23938 36206 23950 36258
rect 21982 36194 22034 36206
rect 28030 36194 28082 36206
rect 28478 36258 28530 36270
rect 28478 36194 28530 36206
rect 29262 36258 29314 36270
rect 29262 36194 29314 36206
rect 34078 36258 34130 36270
rect 34078 36194 34130 36206
rect 37550 36258 37602 36270
rect 37550 36194 37602 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 2494 35922 2546 35934
rect 2494 35858 2546 35870
rect 2606 35922 2658 35934
rect 2606 35858 2658 35870
rect 2830 35922 2882 35934
rect 2830 35858 2882 35870
rect 3502 35922 3554 35934
rect 3502 35858 3554 35870
rect 4622 35922 4674 35934
rect 4622 35858 4674 35870
rect 5742 35922 5794 35934
rect 5742 35858 5794 35870
rect 7646 35922 7698 35934
rect 7646 35858 7698 35870
rect 9998 35922 10050 35934
rect 9998 35858 10050 35870
rect 10222 35922 10274 35934
rect 10222 35858 10274 35870
rect 10334 35922 10386 35934
rect 10334 35858 10386 35870
rect 10670 35922 10722 35934
rect 10670 35858 10722 35870
rect 11790 35922 11842 35934
rect 11790 35858 11842 35870
rect 12014 35922 12066 35934
rect 12014 35858 12066 35870
rect 12574 35922 12626 35934
rect 12574 35858 12626 35870
rect 15038 35922 15090 35934
rect 19742 35922 19794 35934
rect 28702 35922 28754 35934
rect 18722 35870 18734 35922
rect 18786 35870 18798 35922
rect 20850 35870 20862 35922
rect 20914 35870 20926 35922
rect 15038 35858 15090 35870
rect 19742 35858 19794 35870
rect 28702 35858 28754 35870
rect 29150 35922 29202 35934
rect 29150 35858 29202 35870
rect 34750 35922 34802 35934
rect 39342 35922 39394 35934
rect 37650 35870 37662 35922
rect 37714 35870 37726 35922
rect 34750 35858 34802 35870
rect 39342 35858 39394 35870
rect 2270 35810 2322 35822
rect 2270 35746 2322 35758
rect 3726 35810 3778 35822
rect 3726 35746 3778 35758
rect 14814 35810 14866 35822
rect 19966 35810 20018 35822
rect 35646 35810 35698 35822
rect 17714 35758 17726 35810
rect 17778 35758 17790 35810
rect 19170 35758 19182 35810
rect 19234 35758 19246 35810
rect 20514 35758 20526 35810
rect 20578 35758 20590 35810
rect 22866 35758 22878 35810
rect 22930 35758 22942 35810
rect 23874 35758 23886 35810
rect 23938 35758 23950 35810
rect 25442 35758 25454 35810
rect 25506 35758 25518 35810
rect 27458 35758 27470 35810
rect 27522 35758 27534 35810
rect 37762 35758 37774 35810
rect 37826 35758 37838 35810
rect 14814 35746 14866 35758
rect 19966 35746 20018 35758
rect 35646 35746 35698 35758
rect 2718 35698 2770 35710
rect 9662 35698 9714 35710
rect 3266 35646 3278 35698
rect 3330 35646 3342 35698
rect 2718 35634 2770 35646
rect 9662 35634 9714 35646
rect 12126 35698 12178 35710
rect 14702 35698 14754 35710
rect 18734 35698 18786 35710
rect 13906 35646 13918 35698
rect 13970 35646 13982 35698
rect 17602 35646 17614 35698
rect 17666 35646 17678 35698
rect 12126 35634 12178 35646
rect 14702 35634 14754 35646
rect 18734 35634 18786 35646
rect 20078 35698 20130 35710
rect 27806 35698 27858 35710
rect 20962 35646 20974 35698
rect 21026 35646 21038 35698
rect 22978 35646 22990 35698
rect 23042 35646 23054 35698
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 25218 35646 25230 35698
rect 25282 35646 25294 35698
rect 20078 35634 20130 35646
rect 27806 35634 27858 35646
rect 28254 35698 28306 35710
rect 34750 35698 34802 35710
rect 33058 35646 33070 35698
rect 33122 35646 33134 35698
rect 38098 35646 38110 35698
rect 38162 35646 38174 35698
rect 28254 35634 28306 35646
rect 34750 35634 34802 35646
rect 6302 35586 6354 35598
rect 11566 35586 11618 35598
rect 8082 35534 8094 35586
rect 8146 35534 8158 35586
rect 6302 35522 6354 35534
rect 11566 35522 11618 35534
rect 13022 35586 13074 35598
rect 13022 35522 13074 35534
rect 14366 35586 14418 35598
rect 14366 35522 14418 35534
rect 15374 35586 15426 35598
rect 26686 35586 26738 35598
rect 23202 35534 23214 35586
rect 23266 35534 23278 35586
rect 25330 35534 25342 35586
rect 25394 35534 25406 35586
rect 15374 35522 15426 35534
rect 26686 35522 26738 35534
rect 27134 35586 27186 35598
rect 36430 35586 36482 35598
rect 34178 35534 34190 35586
rect 34242 35534 34254 35586
rect 39778 35534 39790 35586
rect 39842 35534 39854 35586
rect 27134 35522 27186 35534
rect 36430 35522 36482 35534
rect 3838 35474 3890 35486
rect 3838 35410 3890 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 12350 35138 12402 35150
rect 11554 35086 11566 35138
rect 11618 35086 11630 35138
rect 12350 35074 12402 35086
rect 18734 35026 18786 35038
rect 2818 34974 2830 35026
rect 2882 34974 2894 35026
rect 9986 34974 9998 35026
rect 10050 34974 10062 35026
rect 14802 34974 14814 35026
rect 14866 34974 14878 35026
rect 17042 34974 17054 35026
rect 17106 34974 17118 35026
rect 18734 34962 18786 34974
rect 26798 35026 26850 35038
rect 41906 34974 41918 35026
rect 41970 34974 41982 35026
rect 26798 34962 26850 34974
rect 2718 34914 2770 34926
rect 2718 34850 2770 34862
rect 6190 34914 6242 34926
rect 8094 34914 8146 34926
rect 6514 34862 6526 34914
rect 6578 34862 6590 34914
rect 6190 34850 6242 34862
rect 8094 34850 8146 34862
rect 8654 34914 8706 34926
rect 8654 34850 8706 34862
rect 10446 34914 10498 34926
rect 10446 34850 10498 34862
rect 10894 34914 10946 34926
rect 12574 34914 12626 34926
rect 19294 34914 19346 34926
rect 12226 34862 12238 34914
rect 12290 34862 12302 34914
rect 13458 34862 13470 34914
rect 13522 34862 13534 34914
rect 14690 34862 14702 34914
rect 14754 34862 14766 34914
rect 16482 34862 16494 34914
rect 16546 34862 16558 34914
rect 16930 34862 16942 34914
rect 16994 34862 17006 34914
rect 10894 34850 10946 34862
rect 12574 34850 12626 34862
rect 19294 34850 19346 34862
rect 19406 34914 19458 34926
rect 19406 34850 19458 34862
rect 20190 34914 20242 34926
rect 20190 34850 20242 34862
rect 20414 34914 20466 34926
rect 26574 34914 26626 34926
rect 20738 34862 20750 34914
rect 20802 34862 20814 34914
rect 22530 34862 22542 34914
rect 22594 34862 22606 34914
rect 23762 34862 23774 34914
rect 23826 34862 23838 34914
rect 25218 34862 25230 34914
rect 25282 34862 25294 34914
rect 20414 34850 20466 34862
rect 26574 34850 26626 34862
rect 27134 34914 27186 34926
rect 27134 34850 27186 34862
rect 27582 34914 27634 34926
rect 27582 34850 27634 34862
rect 27806 34914 27858 34926
rect 27806 34850 27858 34862
rect 28254 34914 28306 34926
rect 28254 34850 28306 34862
rect 29038 34914 29090 34926
rect 29038 34850 29090 34862
rect 32398 34914 32450 34926
rect 32398 34850 32450 34862
rect 32734 34914 32786 34926
rect 35074 34862 35086 34914
rect 35138 34862 35150 34914
rect 36194 34862 36206 34914
rect 36258 34862 36270 34914
rect 37314 34862 37326 34914
rect 37378 34862 37390 34914
rect 39330 34862 39342 34914
rect 39394 34862 39406 34914
rect 32734 34850 32786 34862
rect 2270 34802 2322 34814
rect 2270 34738 2322 34750
rect 2494 34802 2546 34814
rect 2494 34738 2546 34750
rect 2830 34802 2882 34814
rect 2830 34738 2882 34750
rect 5630 34802 5682 34814
rect 11006 34802 11058 34814
rect 7634 34750 7646 34802
rect 7698 34750 7710 34802
rect 5630 34738 5682 34750
rect 11006 34738 11058 34750
rect 11118 34802 11170 34814
rect 11118 34738 11170 34750
rect 13694 34802 13746 34814
rect 18846 34802 18898 34814
rect 27022 34802 27074 34814
rect 14914 34750 14926 34802
rect 14978 34750 14990 34802
rect 15810 34750 15822 34802
rect 15874 34750 15886 34802
rect 16818 34750 16830 34802
rect 16882 34750 16894 34802
rect 21634 34750 21646 34802
rect 21698 34750 21710 34802
rect 23538 34750 23550 34802
rect 23602 34750 23614 34802
rect 25330 34750 25342 34802
rect 25394 34750 25406 34802
rect 25890 34750 25902 34802
rect 25954 34750 25966 34802
rect 13694 34738 13746 34750
rect 18846 34738 18898 34750
rect 27022 34738 27074 34750
rect 29374 34802 29426 34814
rect 29374 34738 29426 34750
rect 29822 34802 29874 34814
rect 29822 34738 29874 34750
rect 33182 34802 33234 34814
rect 39902 34802 39954 34814
rect 34514 34750 34526 34802
rect 34578 34750 34590 34802
rect 36082 34750 36094 34802
rect 36146 34750 36158 34802
rect 37426 34750 37438 34802
rect 37490 34750 37502 34802
rect 33182 34738 33234 34750
rect 39902 34738 39954 34750
rect 12014 34690 12066 34702
rect 12014 34626 12066 34638
rect 12910 34690 12962 34702
rect 12910 34626 12962 34638
rect 19070 34690 19122 34702
rect 19070 34626 19122 34638
rect 20302 34690 20354 34702
rect 27694 34690 27746 34702
rect 22754 34638 22766 34690
rect 22818 34638 22830 34690
rect 26226 34638 26238 34690
rect 26290 34638 26302 34690
rect 20302 34626 20354 34638
rect 27694 34626 27746 34638
rect 28702 34690 28754 34702
rect 28702 34626 28754 34638
rect 29262 34690 29314 34702
rect 29262 34626 29314 34638
rect 30158 34690 30210 34702
rect 30158 34626 30210 34638
rect 30942 34690 30994 34702
rect 30942 34626 30994 34638
rect 31838 34690 31890 34702
rect 41470 34690 41522 34702
rect 34626 34638 34638 34690
rect 34690 34638 34702 34690
rect 37538 34638 37550 34690
rect 37602 34638 37614 34690
rect 31838 34626 31890 34638
rect 41470 34626 41522 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 1710 34354 1762 34366
rect 1710 34290 1762 34302
rect 2494 34354 2546 34366
rect 2494 34290 2546 34302
rect 3950 34354 4002 34366
rect 3950 34290 4002 34302
rect 5406 34354 5458 34366
rect 5406 34290 5458 34302
rect 7870 34354 7922 34366
rect 7870 34290 7922 34302
rect 11566 34354 11618 34366
rect 17278 34354 17330 34366
rect 13906 34302 13918 34354
rect 13970 34302 13982 34354
rect 15810 34302 15822 34354
rect 15874 34302 15886 34354
rect 11566 34290 11618 34302
rect 17278 34290 17330 34302
rect 18062 34354 18114 34366
rect 18062 34290 18114 34302
rect 18510 34354 18562 34366
rect 39230 34354 39282 34366
rect 20066 34302 20078 34354
rect 20130 34302 20142 34354
rect 18510 34290 18562 34302
rect 39230 34290 39282 34302
rect 10558 34242 10610 34254
rect 2034 34190 2046 34242
rect 2098 34190 2110 34242
rect 10558 34178 10610 34190
rect 13134 34242 13186 34254
rect 15934 34242 15986 34254
rect 14354 34190 14366 34242
rect 14418 34190 14430 34242
rect 14802 34190 14814 34242
rect 14866 34190 14878 34242
rect 13134 34178 13186 34190
rect 15934 34178 15986 34190
rect 17502 34242 17554 34254
rect 24222 34242 24274 34254
rect 28030 34242 28082 34254
rect 19842 34190 19854 34242
rect 19906 34190 19918 34242
rect 21858 34190 21870 34242
rect 21922 34190 21934 34242
rect 23874 34190 23886 34242
rect 23938 34190 23950 34242
rect 25890 34190 25902 34242
rect 25954 34190 25966 34242
rect 17502 34178 17554 34190
rect 24222 34178 24274 34190
rect 28030 34178 28082 34190
rect 28142 34242 28194 34254
rect 28142 34178 28194 34190
rect 28254 34242 28306 34254
rect 33954 34190 33966 34242
rect 34018 34190 34030 34242
rect 34850 34190 34862 34242
rect 34914 34190 34926 34242
rect 37762 34190 37774 34242
rect 37826 34190 37838 34242
rect 28254 34178 28306 34190
rect 8542 34130 8594 34142
rect 10670 34130 10722 34142
rect 9650 34078 9662 34130
rect 9714 34078 9726 34130
rect 8542 34066 8594 34078
rect 10670 34066 10722 34078
rect 12462 34130 12514 34142
rect 16718 34130 16770 34142
rect 12898 34078 12910 34130
rect 12962 34078 12974 34130
rect 14130 34078 14142 34130
rect 14194 34078 14206 34130
rect 15250 34078 15262 34130
rect 15314 34078 15326 34130
rect 16146 34078 16158 34130
rect 16210 34078 16222 34130
rect 12462 34066 12514 34078
rect 16718 34066 16770 34078
rect 17614 34130 17666 34142
rect 17614 34066 17666 34078
rect 18398 34130 18450 34142
rect 18398 34066 18450 34078
rect 18622 34130 18674 34142
rect 18622 34066 18674 34078
rect 19070 34130 19122 34142
rect 22206 34130 22258 34142
rect 30830 34130 30882 34142
rect 20402 34078 20414 34130
rect 20466 34078 20478 34130
rect 20962 34078 20974 34130
rect 21026 34078 21038 34130
rect 21186 34078 21198 34130
rect 21250 34078 21262 34130
rect 22642 34078 22654 34130
rect 22706 34078 22718 34130
rect 23538 34078 23550 34130
rect 23602 34078 23614 34130
rect 23986 34078 23998 34130
rect 24050 34078 24062 34130
rect 25330 34078 25342 34130
rect 25394 34078 25406 34130
rect 25554 34078 25566 34130
rect 25618 34078 25630 34130
rect 26226 34078 26238 34130
rect 26290 34078 26302 34130
rect 30370 34078 30382 34130
rect 30434 34078 30446 34130
rect 19070 34066 19122 34078
rect 22206 34066 22258 34078
rect 30830 34066 30882 34078
rect 31390 34130 31442 34142
rect 36654 34130 36706 34142
rect 32498 34078 32510 34130
rect 32562 34078 32574 34130
rect 34402 34078 34414 34130
rect 34466 34078 34478 34130
rect 34738 34078 34750 34130
rect 34802 34078 34814 34130
rect 37090 34078 37102 34130
rect 37154 34078 37166 34130
rect 38658 34078 38670 34130
rect 38722 34078 38734 34130
rect 31390 34066 31442 34078
rect 36654 34066 36706 34078
rect 6638 34018 6690 34030
rect 3490 33966 3502 34018
rect 3554 33966 3566 34018
rect 5842 33966 5854 34018
rect 5906 33966 5918 34018
rect 6638 33954 6690 33966
rect 7086 34018 7138 34030
rect 8318 34018 8370 34030
rect 7410 33966 7422 34018
rect 7474 33966 7486 34018
rect 7086 33954 7138 33966
rect 8318 33954 8370 33966
rect 10110 34018 10162 34030
rect 10110 33954 10162 33966
rect 11118 34018 11170 34030
rect 19518 34018 19570 34030
rect 12002 33966 12014 34018
rect 12066 33966 12078 34018
rect 19058 33966 19070 34018
rect 19122 33966 19134 34018
rect 11118 33954 11170 33966
rect 8878 33906 8930 33918
rect 8878 33842 8930 33854
rect 10558 33906 10610 33918
rect 10994 33854 11006 33906
rect 11058 33903 11070 33906
rect 11666 33903 11678 33906
rect 11058 33857 11678 33903
rect 11058 33854 11070 33857
rect 11666 33854 11678 33857
rect 11730 33854 11742 33906
rect 19073 33903 19119 33966
rect 19518 33954 19570 33966
rect 24670 34018 24722 34030
rect 24670 33954 24722 33966
rect 27246 34018 27298 34030
rect 27246 33954 27298 33966
rect 28814 34018 28866 34030
rect 28814 33954 28866 33966
rect 29262 34018 29314 34030
rect 29262 33954 29314 33966
rect 29934 34018 29986 34030
rect 39790 34018 39842 34030
rect 33618 33966 33630 34018
rect 33682 33966 33694 34018
rect 29934 33954 29986 33966
rect 39790 33954 39842 33966
rect 32398 33906 32450 33918
rect 19618 33903 19630 33906
rect 19073 33857 19630 33903
rect 19618 33854 19630 33857
rect 19682 33854 19694 33906
rect 27570 33854 27582 33906
rect 27634 33854 27646 33906
rect 10558 33842 10610 33854
rect 32398 33842 32450 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 18958 33570 19010 33582
rect 13458 33518 13470 33570
rect 13522 33567 13534 33570
rect 13906 33567 13918 33570
rect 13522 33521 13918 33567
rect 13522 33518 13534 33521
rect 13906 33518 13918 33521
rect 13970 33518 13982 33570
rect 14130 33567 14142 33570
rect 14033 33521 14142 33567
rect 10110 33458 10162 33470
rect 14033 33458 14079 33521
rect 14130 33518 14142 33521
rect 14194 33567 14206 33570
rect 15026 33567 15038 33570
rect 14194 33521 15038 33567
rect 14194 33518 14206 33521
rect 15026 33518 15038 33521
rect 15090 33518 15102 33570
rect 18958 33506 19010 33518
rect 26798 33570 26850 33582
rect 26798 33506 26850 33518
rect 15038 33458 15090 33470
rect 8306 33406 8318 33458
rect 8370 33406 8382 33458
rect 14018 33406 14030 33458
rect 14082 33406 14094 33458
rect 10110 33394 10162 33406
rect 15038 33394 15090 33406
rect 15486 33458 15538 33470
rect 20302 33458 20354 33470
rect 17154 33406 17166 33458
rect 17218 33406 17230 33458
rect 15486 33394 15538 33406
rect 20302 33394 20354 33406
rect 20750 33458 20802 33470
rect 20750 33394 20802 33406
rect 23214 33458 23266 33470
rect 23214 33394 23266 33406
rect 27918 33458 27970 33470
rect 33506 33406 33518 33458
rect 33570 33406 33582 33458
rect 27918 33394 27970 33406
rect 4062 33346 4114 33358
rect 4622 33346 4674 33358
rect 9662 33346 9714 33358
rect 21534 33346 21586 33358
rect 3266 33294 3278 33346
rect 3330 33294 3342 33346
rect 4274 33294 4286 33346
rect 4338 33294 4350 33346
rect 5058 33294 5070 33346
rect 5122 33294 5134 33346
rect 5954 33294 5966 33346
rect 6018 33294 6030 33346
rect 9202 33294 9214 33346
rect 9266 33294 9278 33346
rect 17602 33294 17614 33346
rect 17666 33294 17678 33346
rect 18498 33294 18510 33346
rect 18562 33294 18574 33346
rect 4062 33282 4114 33294
rect 4622 33282 4674 33294
rect 9662 33282 9714 33294
rect 21534 33282 21586 33294
rect 23326 33346 23378 33358
rect 23326 33282 23378 33294
rect 23774 33346 23826 33358
rect 27806 33346 27858 33358
rect 25554 33294 25566 33346
rect 25618 33294 25630 33346
rect 23774 33282 23826 33294
rect 27806 33282 27858 33294
rect 28030 33346 28082 33358
rect 28030 33282 28082 33294
rect 30382 33346 30434 33358
rect 37102 33346 37154 33358
rect 32610 33294 32622 33346
rect 32674 33294 32686 33346
rect 34738 33294 34750 33346
rect 34802 33294 34814 33346
rect 35858 33294 35870 33346
rect 35922 33294 35934 33346
rect 30382 33282 30434 33294
rect 37102 33282 37154 33294
rect 39230 33346 39282 33358
rect 39554 33294 39566 33346
rect 39618 33294 39630 33346
rect 39230 33282 39282 33294
rect 1710 33234 1762 33246
rect 1710 33170 1762 33182
rect 2494 33234 2546 33246
rect 2494 33170 2546 33182
rect 2830 33234 2882 33246
rect 2830 33170 2882 33182
rect 3726 33234 3778 33246
rect 3726 33170 3778 33182
rect 4510 33234 4562 33246
rect 12126 33234 12178 33246
rect 7410 33182 7422 33234
rect 7474 33182 7486 33234
rect 8418 33182 8430 33234
rect 8482 33182 8494 33234
rect 4510 33170 4562 33182
rect 12126 33170 12178 33182
rect 12910 33234 12962 33246
rect 19070 33234 19122 33246
rect 17154 33182 17166 33234
rect 17218 33182 17230 33234
rect 12910 33170 12962 33182
rect 19070 33170 19122 33182
rect 21982 33234 22034 33246
rect 28254 33234 28306 33246
rect 25106 33182 25118 33234
rect 25170 33182 25182 33234
rect 26338 33182 26350 33234
rect 26402 33182 26414 33234
rect 21982 33170 22034 33182
rect 28254 33170 28306 33182
rect 29262 33234 29314 33246
rect 38670 33234 38722 33246
rect 34850 33182 34862 33234
rect 34914 33182 34926 33234
rect 36306 33182 36318 33234
rect 36370 33182 36382 33234
rect 29262 33170 29314 33182
rect 38670 33170 38722 33182
rect 40126 33234 40178 33246
rect 40126 33170 40178 33182
rect 2046 33122 2098 33134
rect 2046 33058 2098 33070
rect 3838 33122 3890 33134
rect 3838 33058 3890 33070
rect 12574 33122 12626 33134
rect 12574 33058 12626 33070
rect 13694 33122 13746 33134
rect 13694 33058 13746 33070
rect 14142 33122 14194 33134
rect 14142 33058 14194 33070
rect 14590 33122 14642 33134
rect 14590 33058 14642 33070
rect 16382 33122 16434 33134
rect 16382 33058 16434 33070
rect 18286 33122 18338 33134
rect 18286 33058 18338 33070
rect 18958 33122 19010 33134
rect 18958 33058 19010 33070
rect 19518 33122 19570 33134
rect 19518 33058 19570 33070
rect 22430 33122 22482 33134
rect 22430 33058 22482 33070
rect 22878 33122 22930 33134
rect 22878 33058 22930 33070
rect 23102 33122 23154 33134
rect 23102 33058 23154 33070
rect 27694 33122 27746 33134
rect 27694 33058 27746 33070
rect 30942 33122 30994 33134
rect 37214 33122 37266 33134
rect 35298 33070 35310 33122
rect 35362 33070 35374 33122
rect 38994 33070 39006 33122
rect 39058 33070 39070 33122
rect 30942 33058 30994 33070
rect 37214 33058 37266 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 19182 32786 19234 32798
rect 5170 32734 5182 32786
rect 5234 32734 5246 32786
rect 13458 32734 13470 32786
rect 13522 32734 13534 32786
rect 19182 32722 19234 32734
rect 24670 32786 24722 32798
rect 24670 32722 24722 32734
rect 28926 32786 28978 32798
rect 28926 32722 28978 32734
rect 14030 32674 14082 32686
rect 5394 32622 5406 32674
rect 5458 32622 5470 32674
rect 14030 32610 14082 32622
rect 14366 32674 14418 32686
rect 14366 32610 14418 32622
rect 16830 32674 16882 32686
rect 28366 32674 28418 32686
rect 17938 32622 17950 32674
rect 18002 32622 18014 32674
rect 21858 32622 21870 32674
rect 21922 32622 21934 32674
rect 22306 32622 22318 32674
rect 22370 32622 22382 32674
rect 16830 32610 16882 32622
rect 28366 32610 28418 32622
rect 28478 32674 28530 32686
rect 28478 32610 28530 32622
rect 33630 32674 33682 32686
rect 33630 32610 33682 32622
rect 36206 32674 36258 32686
rect 36206 32610 36258 32622
rect 7310 32562 7362 32574
rect 2370 32510 2382 32562
rect 2434 32510 2446 32562
rect 3266 32510 3278 32562
rect 3330 32510 3342 32562
rect 3602 32510 3614 32562
rect 3666 32510 3678 32562
rect 4946 32510 4958 32562
rect 5010 32510 5022 32562
rect 6514 32510 6526 32562
rect 6578 32510 6590 32562
rect 7310 32498 7362 32510
rect 8990 32562 9042 32574
rect 28142 32562 28194 32574
rect 10322 32510 10334 32562
rect 10386 32510 10398 32562
rect 12114 32510 12126 32562
rect 12178 32510 12190 32562
rect 13234 32510 13246 32562
rect 13298 32510 13310 32562
rect 17714 32510 17726 32562
rect 17778 32510 17790 32562
rect 18834 32510 18846 32562
rect 18898 32510 18910 32562
rect 21634 32510 21646 32562
rect 21698 32510 21710 32562
rect 23650 32510 23662 32562
rect 23714 32510 23726 32562
rect 25330 32510 25342 32562
rect 25394 32510 25406 32562
rect 26338 32510 26350 32562
rect 26402 32510 26414 32562
rect 27458 32510 27470 32562
rect 27522 32510 27534 32562
rect 33058 32510 33070 32562
rect 33122 32510 33134 32562
rect 35074 32510 35086 32562
rect 35138 32510 35150 32562
rect 38434 32510 38446 32562
rect 38498 32510 38510 32562
rect 40002 32510 40014 32562
rect 40066 32510 40078 32562
rect 8990 32498 9042 32510
rect 28142 32498 28194 32510
rect 15486 32450 15538 32462
rect 8530 32398 8542 32450
rect 8594 32398 8606 32450
rect 10658 32398 10670 32450
rect 10722 32398 10734 32450
rect 12450 32398 12462 32450
rect 12514 32398 12526 32450
rect 14802 32398 14814 32450
rect 14866 32398 14878 32450
rect 15486 32386 15538 32398
rect 16494 32450 16546 32462
rect 21422 32450 21474 32462
rect 34862 32450 34914 32462
rect 18162 32398 18174 32450
rect 18226 32398 18238 32450
rect 23202 32398 23214 32450
rect 23266 32398 23278 32450
rect 37538 32398 37550 32450
rect 37602 32398 37614 32450
rect 39554 32398 39566 32450
rect 39618 32398 39630 32450
rect 16494 32386 16546 32398
rect 21422 32386 21474 32398
rect 34862 32386 34914 32398
rect 26786 32286 26798 32338
rect 26850 32286 26862 32338
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 17390 32002 17442 32014
rect 17390 31938 17442 31950
rect 20414 31890 20466 31902
rect 27134 31890 27186 31902
rect 2594 31838 2606 31890
rect 2658 31838 2670 31890
rect 3490 31838 3502 31890
rect 3554 31838 3566 31890
rect 18274 31838 18286 31890
rect 18338 31838 18350 31890
rect 24546 31838 24558 31890
rect 24610 31838 24622 31890
rect 20414 31826 20466 31838
rect 27134 31826 27186 31838
rect 29150 31890 29202 31902
rect 30482 31838 30494 31890
rect 30546 31838 30558 31890
rect 29150 31826 29202 31838
rect 3054 31778 3106 31790
rect 13470 31778 13522 31790
rect 8978 31726 8990 31778
rect 9042 31726 9054 31778
rect 9314 31726 9326 31778
rect 9378 31726 9390 31778
rect 9650 31726 9662 31778
rect 9714 31726 9726 31778
rect 10994 31726 11006 31778
rect 11058 31726 11070 31778
rect 12786 31726 12798 31778
rect 12850 31726 12862 31778
rect 3054 31714 3106 31726
rect 13470 31714 13522 31726
rect 14030 31778 14082 31790
rect 19854 31778 19906 31790
rect 15250 31726 15262 31778
rect 15314 31726 15326 31778
rect 15810 31726 15822 31778
rect 15874 31726 15886 31778
rect 16594 31726 16606 31778
rect 16658 31726 16670 31778
rect 17042 31726 17054 31778
rect 17106 31726 17118 31778
rect 17714 31726 17726 31778
rect 17778 31726 17790 31778
rect 18498 31726 18510 31778
rect 18562 31726 18574 31778
rect 14030 31714 14082 31726
rect 19854 31714 19906 31726
rect 20190 31778 20242 31790
rect 20190 31714 20242 31726
rect 20750 31778 20802 31790
rect 20750 31714 20802 31726
rect 22430 31778 22482 31790
rect 26798 31778 26850 31790
rect 22866 31726 22878 31778
rect 22930 31726 22942 31778
rect 24882 31726 24894 31778
rect 24946 31726 24958 31778
rect 22430 31714 22482 31726
rect 26798 31714 26850 31726
rect 27358 31778 27410 31790
rect 27358 31714 27410 31726
rect 33966 31778 34018 31790
rect 39118 31778 39170 31790
rect 34290 31726 34302 31778
rect 34354 31726 34366 31778
rect 36978 31726 36990 31778
rect 37042 31726 37054 31778
rect 33966 31714 34018 31726
rect 39118 31714 39170 31726
rect 14590 31666 14642 31678
rect 11442 31614 11454 31666
rect 11506 31614 11518 31666
rect 14590 31602 14642 31614
rect 14814 31666 14866 31678
rect 14814 31602 14866 31614
rect 15038 31666 15090 31678
rect 15038 31602 15090 31614
rect 16046 31666 16098 31678
rect 33406 31666 33458 31678
rect 39678 31666 39730 31678
rect 17938 31614 17950 31666
rect 18002 31614 18014 31666
rect 24210 31614 24222 31666
rect 24274 31614 24286 31666
rect 25218 31614 25230 31666
rect 25282 31614 25294 31666
rect 27794 31614 27806 31666
rect 27858 31614 27870 31666
rect 28018 31614 28030 31666
rect 28082 31614 28094 31666
rect 36082 31614 36094 31666
rect 36146 31614 36158 31666
rect 37090 31614 37102 31666
rect 37154 31614 37166 31666
rect 16046 31602 16098 31614
rect 33406 31602 33458 31614
rect 39678 31602 39730 31614
rect 3950 31554 4002 31566
rect 14926 31554 14978 31566
rect 19630 31554 19682 31566
rect 12898 31502 12910 31554
rect 12962 31502 12974 31554
rect 18946 31502 18958 31554
rect 19010 31502 19022 31554
rect 3950 31490 4002 31502
rect 14926 31490 14978 31502
rect 19630 31490 19682 31502
rect 19742 31554 19794 31566
rect 19742 31490 19794 31502
rect 20302 31554 20354 31566
rect 20302 31490 20354 31502
rect 21422 31554 21474 31566
rect 21422 31490 21474 31502
rect 29710 31554 29762 31566
rect 29710 31490 29762 31502
rect 30942 31554 30994 31566
rect 32386 31502 32398 31554
rect 32450 31502 32462 31554
rect 37202 31502 37214 31554
rect 37266 31502 37278 31554
rect 30942 31490 30994 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 2270 31218 2322 31230
rect 2270 31154 2322 31166
rect 9102 31218 9154 31230
rect 13694 31218 13746 31230
rect 10882 31166 10894 31218
rect 10946 31166 10958 31218
rect 9102 31154 9154 31166
rect 13694 31154 13746 31166
rect 14142 31218 14194 31230
rect 14142 31154 14194 31166
rect 14366 31218 14418 31230
rect 14366 31154 14418 31166
rect 15150 31218 15202 31230
rect 15150 31154 15202 31166
rect 15486 31218 15538 31230
rect 15486 31154 15538 31166
rect 16270 31218 16322 31230
rect 16270 31154 16322 31166
rect 17838 31218 17890 31230
rect 17838 31154 17890 31166
rect 19070 31218 19122 31230
rect 19070 31154 19122 31166
rect 20974 31218 21026 31230
rect 20974 31154 21026 31166
rect 24222 31218 24274 31230
rect 24222 31154 24274 31166
rect 24782 31218 24834 31230
rect 24782 31154 24834 31166
rect 25790 31218 25842 31230
rect 25790 31154 25842 31166
rect 26462 31218 26514 31230
rect 26462 31154 26514 31166
rect 26686 31218 26738 31230
rect 26686 31154 26738 31166
rect 27806 31218 27858 31230
rect 27806 31154 27858 31166
rect 28478 31218 28530 31230
rect 28478 31154 28530 31166
rect 28814 31218 28866 31230
rect 28814 31154 28866 31166
rect 29038 31218 29090 31230
rect 33170 31166 33182 31218
rect 33234 31166 33246 31218
rect 29038 31154 29090 31166
rect 13918 31106 13970 31118
rect 3042 31054 3054 31106
rect 3106 31054 3118 31106
rect 4386 31054 4398 31106
rect 4450 31054 4462 31106
rect 5618 31054 5630 31106
rect 5682 31054 5694 31106
rect 12338 31054 12350 31106
rect 12402 31054 12414 31106
rect 13918 31042 13970 31054
rect 17390 31106 17442 31118
rect 17390 31042 17442 31054
rect 17614 31106 17666 31118
rect 17614 31042 17666 31054
rect 18062 31106 18114 31118
rect 18062 31042 18114 31054
rect 20078 31106 20130 31118
rect 20078 31042 20130 31054
rect 20302 31106 20354 31118
rect 20302 31042 20354 31054
rect 34302 31106 34354 31118
rect 34302 31042 34354 31054
rect 35758 31106 35810 31118
rect 35758 31042 35810 31054
rect 6974 30994 7026 31006
rect 16158 30994 16210 31006
rect 2146 30942 2158 30994
rect 2210 30942 2222 30994
rect 3490 30942 3502 30994
rect 3554 30942 3566 30994
rect 4274 30942 4286 30994
rect 4338 30942 4350 30994
rect 10098 30942 10110 30994
rect 10162 30942 10174 30994
rect 10994 30942 11006 30994
rect 11058 30942 11070 30994
rect 11890 30942 11902 30994
rect 11954 30942 11966 30994
rect 14578 30942 14590 30994
rect 14642 30942 14654 30994
rect 6974 30930 7026 30942
rect 16158 30930 16210 30942
rect 18622 30994 18674 31006
rect 18622 30930 18674 30942
rect 18734 30994 18786 31006
rect 18734 30930 18786 30942
rect 18958 30994 19010 31006
rect 18958 30930 19010 30942
rect 20638 30994 20690 31006
rect 20638 30930 20690 30942
rect 26014 30994 26066 31006
rect 26014 30930 26066 30942
rect 27246 30994 27298 31006
rect 27246 30930 27298 30942
rect 27694 30994 27746 31006
rect 27694 30930 27746 30942
rect 27918 30994 27970 31006
rect 27918 30930 27970 30942
rect 29486 30994 29538 31006
rect 34850 30942 34862 30994
rect 34914 30942 34926 30994
rect 36866 30942 36878 30994
rect 36930 30942 36942 30994
rect 38210 30942 38222 30994
rect 38274 30942 38286 30994
rect 29486 30930 29538 30942
rect 7534 30882 7586 30894
rect 3378 30830 3390 30882
rect 3442 30830 3454 30882
rect 6290 30830 6302 30882
rect 6354 30830 6366 30882
rect 7534 30818 7586 30830
rect 8654 30882 8706 30894
rect 8654 30818 8706 30830
rect 14254 30882 14306 30894
rect 14254 30818 14306 30830
rect 16830 30882 16882 30894
rect 16830 30818 16882 30830
rect 18174 30882 18226 30894
rect 18174 30818 18226 30830
rect 18846 30882 18898 30894
rect 18846 30818 18898 30830
rect 19630 30882 19682 30894
rect 19630 30818 19682 30830
rect 21422 30882 21474 30894
rect 21422 30818 21474 30830
rect 21870 30882 21922 30894
rect 26574 30882 26626 30894
rect 25330 30830 25342 30882
rect 25394 30830 25406 30882
rect 21870 30818 21922 30830
rect 26574 30818 26626 30830
rect 28926 30882 28978 30894
rect 37314 30830 37326 30882
rect 37378 30830 37390 30882
rect 28926 30818 28978 30830
rect 16270 30770 16322 30782
rect 8642 30718 8654 30770
rect 8706 30767 8718 30770
rect 9090 30767 9102 30770
rect 8706 30721 9102 30767
rect 8706 30718 8718 30721
rect 9090 30718 9102 30721
rect 9154 30718 9166 30770
rect 15138 30718 15150 30770
rect 15202 30767 15214 30770
rect 15698 30767 15710 30770
rect 15202 30721 15710 30767
rect 15202 30718 15214 30721
rect 15698 30718 15710 30721
rect 15762 30718 15774 30770
rect 16270 30706 16322 30718
rect 20862 30770 20914 30782
rect 20862 30706 20914 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 21870 30434 21922 30446
rect 14354 30382 14366 30434
rect 14418 30431 14430 30434
rect 14914 30431 14926 30434
rect 14418 30385 14926 30431
rect 14418 30382 14430 30385
rect 14914 30382 14926 30385
rect 14978 30382 14990 30434
rect 21870 30370 21922 30382
rect 26014 30434 26066 30446
rect 26014 30370 26066 30382
rect 6526 30322 6578 30334
rect 11790 30322 11842 30334
rect 9202 30270 9214 30322
rect 9266 30270 9278 30322
rect 6526 30258 6578 30270
rect 11790 30258 11842 30270
rect 14926 30322 14978 30334
rect 14926 30258 14978 30270
rect 27022 30322 27074 30334
rect 34414 30322 34466 30334
rect 30482 30270 30494 30322
rect 30546 30270 30558 30322
rect 27022 30258 27074 30270
rect 34414 30258 34466 30270
rect 36206 30322 36258 30334
rect 36206 30258 36258 30270
rect 1710 30210 1762 30222
rect 1710 30146 1762 30158
rect 4734 30210 4786 30222
rect 6414 30210 6466 30222
rect 9102 30210 9154 30222
rect 6178 30158 6190 30210
rect 6242 30158 6254 30210
rect 6850 30158 6862 30210
rect 6914 30158 6926 30210
rect 7858 30158 7870 30210
rect 7922 30158 7934 30210
rect 8418 30158 8430 30210
rect 8482 30158 8494 30210
rect 4734 30146 4786 30158
rect 6414 30146 6466 30158
rect 9102 30146 9154 30158
rect 9886 30210 9938 30222
rect 9886 30146 9938 30158
rect 12910 30210 12962 30222
rect 14030 30210 14082 30222
rect 13570 30158 13582 30210
rect 13634 30158 13646 30210
rect 12910 30146 12962 30158
rect 14030 30146 14082 30158
rect 15486 30210 15538 30222
rect 15486 30146 15538 30158
rect 17278 30210 17330 30222
rect 17278 30146 17330 30158
rect 17502 30210 17554 30222
rect 21534 30210 21586 30222
rect 18274 30158 18286 30210
rect 18338 30158 18350 30210
rect 19282 30158 19294 30210
rect 19346 30158 19358 30210
rect 19954 30158 19966 30210
rect 20018 30158 20030 30210
rect 17502 30146 17554 30158
rect 21534 30146 21586 30158
rect 21758 30210 21810 30222
rect 23550 30210 23602 30222
rect 22418 30158 22430 30210
rect 22482 30158 22494 30210
rect 21758 30146 21810 30158
rect 23550 30146 23602 30158
rect 25006 30210 25058 30222
rect 25006 30146 25058 30158
rect 25118 30210 25170 30222
rect 28590 30210 28642 30222
rect 31502 30210 31554 30222
rect 25442 30158 25454 30210
rect 25506 30158 25518 30210
rect 26338 30158 26350 30210
rect 26402 30158 26414 30210
rect 26562 30158 26574 30210
rect 26626 30158 26638 30210
rect 30930 30158 30942 30210
rect 30994 30158 31006 30210
rect 31938 30158 31950 30210
rect 32002 30158 32014 30210
rect 34850 30158 34862 30210
rect 34914 30158 34926 30210
rect 35858 30158 35870 30210
rect 35922 30158 35934 30210
rect 25118 30146 25170 30158
rect 28590 30146 28642 30158
rect 31502 30146 31554 30158
rect 2046 30098 2098 30110
rect 2046 30034 2098 30046
rect 2382 30098 2434 30110
rect 2382 30034 2434 30046
rect 4174 30098 4226 30110
rect 4174 30034 4226 30046
rect 5070 30098 5122 30110
rect 11230 30098 11282 30110
rect 7522 30046 7534 30098
rect 7586 30046 7598 30098
rect 9650 30046 9662 30098
rect 9714 30046 9726 30098
rect 5070 30034 5122 30046
rect 11230 30034 11282 30046
rect 11678 30098 11730 30110
rect 11678 30034 11730 30046
rect 12126 30098 12178 30110
rect 12126 30034 12178 30046
rect 12574 30098 12626 30110
rect 12574 30034 12626 30046
rect 12686 30098 12738 30110
rect 12686 30034 12738 30046
rect 20414 30098 20466 30110
rect 20414 30034 20466 30046
rect 21310 30098 21362 30110
rect 21310 30034 21362 30046
rect 21982 30098 22034 30110
rect 23326 30098 23378 30110
rect 25230 30098 25282 30110
rect 22642 30046 22654 30098
rect 22706 30046 22718 30098
rect 23090 30046 23102 30098
rect 23154 30046 23166 30098
rect 23986 30046 23998 30098
rect 24050 30046 24062 30098
rect 24322 30046 24334 30098
rect 24386 30046 24398 30098
rect 21982 30034 22034 30046
rect 23326 30034 23378 30046
rect 25230 30034 25282 30046
rect 25902 30098 25954 30110
rect 25902 30034 25954 30046
rect 28142 30098 28194 30110
rect 28142 30034 28194 30046
rect 2718 29986 2770 29998
rect 2718 29922 2770 29934
rect 3166 29986 3218 29998
rect 3166 29922 3218 29934
rect 4622 29986 4674 29998
rect 4622 29922 4674 29934
rect 4958 29986 5010 29998
rect 4958 29922 5010 29934
rect 5854 29986 5906 29998
rect 5854 29922 5906 29934
rect 6638 29986 6690 29998
rect 6638 29922 6690 29934
rect 10670 29986 10722 29998
rect 10670 29922 10722 29934
rect 11566 29986 11618 29998
rect 11566 29922 11618 29934
rect 11902 29986 11954 29998
rect 11902 29922 11954 29934
rect 14478 29986 14530 29998
rect 14478 29922 14530 29934
rect 26126 29986 26178 29998
rect 26126 29922 26178 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 1822 29650 1874 29662
rect 7086 29650 7138 29662
rect 6178 29598 6190 29650
rect 6242 29598 6254 29650
rect 1822 29586 1874 29598
rect 7086 29586 7138 29598
rect 11678 29650 11730 29662
rect 15710 29650 15762 29662
rect 12674 29598 12686 29650
rect 12738 29598 12750 29650
rect 15138 29598 15150 29650
rect 15202 29598 15214 29650
rect 11678 29586 11730 29598
rect 2818 29486 2830 29538
rect 2882 29486 2894 29538
rect 6402 29486 6414 29538
rect 6466 29486 6478 29538
rect 7522 29486 7534 29538
rect 7586 29486 7598 29538
rect 9762 29486 9774 29538
rect 9826 29486 9838 29538
rect 12462 29426 12514 29438
rect 2258 29374 2270 29426
rect 2322 29374 2334 29426
rect 4610 29374 4622 29426
rect 4674 29374 4686 29426
rect 5730 29374 5742 29426
rect 5794 29374 5806 29426
rect 7970 29374 7982 29426
rect 8034 29374 8046 29426
rect 8866 29374 8878 29426
rect 8930 29374 8942 29426
rect 9650 29374 9662 29426
rect 9714 29374 9726 29426
rect 10210 29374 10222 29426
rect 10274 29374 10286 29426
rect 10994 29374 11006 29426
rect 11058 29374 11070 29426
rect 12462 29362 12514 29374
rect 7646 29314 7698 29326
rect 12002 29262 12014 29314
rect 12066 29262 12078 29314
rect 7646 29250 7698 29262
rect 10222 29202 10274 29214
rect 12689 29202 12735 29598
rect 15710 29586 15762 29598
rect 16158 29650 16210 29662
rect 16158 29586 16210 29598
rect 18958 29650 19010 29662
rect 18958 29586 19010 29598
rect 19518 29650 19570 29662
rect 19518 29586 19570 29598
rect 20078 29650 20130 29662
rect 20078 29586 20130 29598
rect 20862 29650 20914 29662
rect 20862 29586 20914 29598
rect 23438 29650 23490 29662
rect 23438 29586 23490 29598
rect 23774 29650 23826 29662
rect 23774 29586 23826 29598
rect 23998 29650 24050 29662
rect 23998 29586 24050 29598
rect 24222 29650 24274 29662
rect 24222 29586 24274 29598
rect 25566 29650 25618 29662
rect 25566 29586 25618 29598
rect 26014 29650 26066 29662
rect 26014 29586 26066 29598
rect 27246 29650 27298 29662
rect 27246 29586 27298 29598
rect 27806 29650 27858 29662
rect 35634 29598 35646 29650
rect 35698 29598 35710 29650
rect 27806 29586 27858 29598
rect 13694 29538 13746 29550
rect 13694 29474 13746 29486
rect 14702 29538 14754 29550
rect 14702 29474 14754 29486
rect 20414 29538 20466 29550
rect 20414 29474 20466 29486
rect 27582 29538 27634 29550
rect 27582 29474 27634 29486
rect 27918 29538 27970 29550
rect 37326 29538 37378 29550
rect 28578 29486 28590 29538
rect 28642 29486 28654 29538
rect 34178 29486 34190 29538
rect 34242 29486 34254 29538
rect 27918 29474 27970 29486
rect 37326 29474 37378 29486
rect 14590 29426 14642 29438
rect 19966 29426 20018 29438
rect 14354 29374 14366 29426
rect 14418 29374 14430 29426
rect 19730 29374 19742 29426
rect 19794 29374 19806 29426
rect 14590 29362 14642 29374
rect 19966 29362 20018 29374
rect 20190 29426 20242 29438
rect 20190 29362 20242 29374
rect 21198 29426 21250 29438
rect 21198 29362 21250 29374
rect 21758 29426 21810 29438
rect 21758 29362 21810 29374
rect 22206 29426 22258 29438
rect 22206 29362 22258 29374
rect 24334 29426 24386 29438
rect 24334 29362 24386 29374
rect 28030 29426 28082 29438
rect 28030 29362 28082 29374
rect 28366 29426 28418 29438
rect 35870 29426 35922 29438
rect 28914 29374 28926 29426
rect 28978 29374 28990 29426
rect 29586 29374 29598 29426
rect 29650 29374 29662 29426
rect 28366 29362 28418 29374
rect 35870 29362 35922 29374
rect 37886 29426 37938 29438
rect 37886 29362 37938 29374
rect 22654 29314 22706 29326
rect 22654 29250 22706 29262
rect 26686 29314 26738 29326
rect 26686 29250 26738 29262
rect 13134 29202 13186 29214
rect 12674 29150 12686 29202
rect 12738 29150 12750 29202
rect 10222 29138 10274 29150
rect 13134 29138 13186 29150
rect 13358 29202 13410 29214
rect 13358 29138 13410 29150
rect 13806 29202 13858 29214
rect 13806 29138 13858 29150
rect 13918 29202 13970 29214
rect 29934 29202 29986 29214
rect 15362 29150 15374 29202
rect 15426 29199 15438 29202
rect 16146 29199 16158 29202
rect 15426 29153 16158 29199
rect 15426 29150 15438 29153
rect 16146 29150 16158 29153
rect 16210 29150 16222 29202
rect 25778 29150 25790 29202
rect 25842 29199 25854 29202
rect 26114 29199 26126 29202
rect 25842 29153 26126 29199
rect 25842 29150 25854 29153
rect 26114 29150 26126 29153
rect 26178 29150 26190 29202
rect 13918 29138 13970 29150
rect 29934 29138 29986 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 21534 28866 21586 28878
rect 30146 28814 30158 28866
rect 30210 28814 30222 28866
rect 21534 28802 21586 28814
rect 2606 28754 2658 28766
rect 6078 28754 6130 28766
rect 11790 28754 11842 28766
rect 3826 28702 3838 28754
rect 3890 28702 3902 28754
rect 10658 28702 10670 28754
rect 10722 28702 10734 28754
rect 2606 28690 2658 28702
rect 6078 28690 6130 28702
rect 11790 28690 11842 28702
rect 12126 28754 12178 28766
rect 12126 28690 12178 28702
rect 12686 28754 12738 28766
rect 12686 28690 12738 28702
rect 14478 28754 14530 28766
rect 14478 28690 14530 28702
rect 15038 28754 15090 28766
rect 15038 28690 15090 28702
rect 16606 28754 16658 28766
rect 16606 28690 16658 28702
rect 20078 28754 20130 28766
rect 26910 28754 26962 28766
rect 24546 28702 24558 28754
rect 24610 28702 24622 28754
rect 26338 28702 26350 28754
rect 26402 28702 26414 28754
rect 20078 28690 20130 28702
rect 26910 28690 26962 28702
rect 27470 28754 27522 28766
rect 27470 28690 27522 28702
rect 2830 28642 2882 28654
rect 10110 28642 10162 28654
rect 15150 28642 15202 28654
rect 2258 28590 2270 28642
rect 2322 28590 2334 28642
rect 3938 28590 3950 28642
rect 4002 28590 4014 28642
rect 6402 28590 6414 28642
rect 6466 28590 6478 28642
rect 10546 28590 10558 28642
rect 10610 28590 10622 28642
rect 11218 28590 11230 28642
rect 11282 28590 11294 28642
rect 2830 28578 2882 28590
rect 10110 28578 10162 28590
rect 15150 28578 15202 28590
rect 15262 28642 15314 28654
rect 15262 28578 15314 28590
rect 16046 28642 16098 28654
rect 16046 28578 16098 28590
rect 18510 28642 18562 28654
rect 18510 28578 18562 28590
rect 18846 28642 18898 28654
rect 18846 28578 18898 28590
rect 19294 28642 19346 28654
rect 19294 28578 19346 28590
rect 20414 28642 20466 28654
rect 20414 28578 20466 28590
rect 20750 28642 20802 28654
rect 20750 28578 20802 28590
rect 21982 28642 22034 28654
rect 21982 28578 22034 28590
rect 22542 28642 22594 28654
rect 25118 28642 25170 28654
rect 28590 28642 28642 28654
rect 23314 28590 23326 28642
rect 23378 28590 23390 28642
rect 24658 28590 24670 28642
rect 24722 28590 24734 28642
rect 26002 28590 26014 28642
rect 26066 28590 26078 28642
rect 22542 28578 22594 28590
rect 25118 28578 25170 28590
rect 28590 28578 28642 28590
rect 29150 28642 29202 28654
rect 29150 28578 29202 28590
rect 29262 28642 29314 28654
rect 29262 28578 29314 28590
rect 29486 28642 29538 28654
rect 29486 28578 29538 28590
rect 29710 28642 29762 28654
rect 29710 28578 29762 28590
rect 2494 28530 2546 28542
rect 2494 28466 2546 28478
rect 3278 28530 3330 28542
rect 3278 28466 3330 28478
rect 6974 28530 7026 28542
rect 11006 28530 11058 28542
rect 10210 28478 10222 28530
rect 10274 28478 10286 28530
rect 6974 28466 7026 28478
rect 11006 28466 11058 28478
rect 14702 28530 14754 28542
rect 14702 28466 14754 28478
rect 18734 28530 18786 28542
rect 18734 28466 18786 28478
rect 21646 28530 21698 28542
rect 21646 28466 21698 28478
rect 23438 28530 23490 28542
rect 28254 28530 28306 28542
rect 24210 28478 24222 28530
rect 24274 28478 24286 28530
rect 23438 28466 23490 28478
rect 28254 28466 28306 28478
rect 28366 28530 28418 28542
rect 28366 28466 28418 28478
rect 2718 28418 2770 28430
rect 2718 28354 2770 28366
rect 3502 28418 3554 28430
rect 3502 28354 3554 28366
rect 3726 28418 3778 28430
rect 10782 28418 10834 28430
rect 6626 28366 6638 28418
rect 6690 28366 6702 28418
rect 3726 28354 3778 28366
rect 10782 28354 10834 28366
rect 14926 28418 14978 28430
rect 14926 28354 14978 28366
rect 18286 28418 18338 28430
rect 18286 28354 18338 28366
rect 20526 28418 20578 28430
rect 20526 28354 20578 28366
rect 21534 28418 21586 28430
rect 21534 28354 21586 28366
rect 28030 28418 28082 28430
rect 28030 28354 28082 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 2046 28082 2098 28094
rect 2046 28018 2098 28030
rect 4734 28082 4786 28094
rect 4734 28018 4786 28030
rect 5182 28082 5234 28094
rect 5182 28018 5234 28030
rect 7086 28082 7138 28094
rect 8542 28082 8594 28094
rect 7970 28030 7982 28082
rect 8034 28030 8046 28082
rect 7086 28018 7138 28030
rect 8542 28018 8594 28030
rect 8654 28082 8706 28094
rect 8654 28018 8706 28030
rect 8766 28082 8818 28094
rect 8766 28018 8818 28030
rect 11454 28082 11506 28094
rect 16718 28082 16770 28094
rect 13010 28030 13022 28082
rect 13074 28030 13086 28082
rect 16258 28030 16270 28082
rect 16322 28030 16334 28082
rect 11454 28018 11506 28030
rect 16718 28018 16770 28030
rect 18174 28082 18226 28094
rect 18174 28018 18226 28030
rect 22990 28082 23042 28094
rect 22990 28018 23042 28030
rect 25454 28082 25506 28094
rect 25454 28018 25506 28030
rect 25790 28082 25842 28094
rect 29934 28082 29986 28094
rect 27010 28030 27022 28082
rect 27074 28030 27086 28082
rect 25790 28018 25842 28030
rect 29934 28018 29986 28030
rect 30830 28082 30882 28094
rect 30830 28018 30882 28030
rect 4174 27970 4226 27982
rect 4174 27906 4226 27918
rect 4958 27970 5010 27982
rect 4958 27906 5010 27918
rect 5966 27970 6018 27982
rect 5966 27906 6018 27918
rect 8990 27970 9042 27982
rect 18398 27970 18450 27982
rect 21646 27970 21698 27982
rect 30270 27970 30322 27982
rect 12338 27918 12350 27970
rect 12402 27918 12414 27970
rect 19618 27918 19630 27970
rect 19682 27918 19694 27970
rect 20626 27918 20638 27970
rect 20690 27918 20702 27970
rect 20962 27918 20974 27970
rect 21026 27918 21038 27970
rect 27346 27918 27358 27970
rect 27410 27918 27422 27970
rect 8990 27906 9042 27918
rect 18398 27906 18450 27918
rect 21646 27906 21698 27918
rect 30270 27906 30322 27918
rect 1710 27858 1762 27870
rect 1710 27794 1762 27806
rect 5518 27858 5570 27870
rect 8430 27858 8482 27870
rect 15710 27858 15762 27870
rect 5730 27806 5742 27858
rect 5794 27806 5806 27858
rect 6626 27806 6638 27858
rect 6690 27806 6702 27858
rect 6962 27806 6974 27858
rect 7026 27806 7038 27858
rect 7746 27806 7758 27858
rect 7810 27806 7822 27858
rect 10546 27806 10558 27858
rect 10610 27806 10622 27858
rect 12114 27806 12126 27858
rect 12178 27806 12190 27858
rect 13682 27806 13694 27858
rect 13746 27806 13758 27858
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 15474 27806 15486 27858
rect 15538 27806 15550 27858
rect 5518 27794 5570 27806
rect 8430 27794 8482 27806
rect 15710 27794 15762 27806
rect 15822 27858 15874 27870
rect 15822 27794 15874 27806
rect 16606 27858 16658 27870
rect 16606 27794 16658 27806
rect 17726 27858 17778 27870
rect 17726 27794 17778 27806
rect 17950 27858 18002 27870
rect 21534 27858 21586 27870
rect 18722 27806 18734 27858
rect 18786 27806 18798 27858
rect 19394 27806 19406 27858
rect 19458 27806 19470 27858
rect 19954 27806 19966 27858
rect 20018 27806 20030 27858
rect 17950 27794 18002 27806
rect 21534 27794 21586 27806
rect 25678 27858 25730 27870
rect 25678 27794 25730 27806
rect 25902 27858 25954 27870
rect 25902 27794 25954 27806
rect 26462 27858 26514 27870
rect 28142 27858 28194 27870
rect 27570 27806 27582 27858
rect 27634 27806 27646 27858
rect 26462 27794 26514 27806
rect 28142 27794 28194 27806
rect 29374 27858 29426 27870
rect 29374 27794 29426 27806
rect 2494 27746 2546 27758
rect 2494 27682 2546 27694
rect 5294 27746 5346 27758
rect 24670 27746 24722 27758
rect 9986 27694 9998 27746
rect 10050 27694 10062 27746
rect 5294 27682 5346 27694
rect 24670 27682 24722 27694
rect 16718 27634 16770 27646
rect 16718 27570 16770 27582
rect 17838 27634 17890 27646
rect 17838 27570 17890 27582
rect 26686 27634 26738 27646
rect 26686 27570 26738 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 17602 27246 17614 27298
rect 17666 27295 17678 27298
rect 17826 27295 17838 27298
rect 17666 27249 17838 27295
rect 17666 27246 17678 27249
rect 17826 27246 17838 27249
rect 17890 27246 17902 27298
rect 24658 27246 24670 27298
rect 24722 27246 24734 27298
rect 4622 27186 4674 27198
rect 3714 27134 3726 27186
rect 3778 27134 3790 27186
rect 4622 27122 4674 27134
rect 6414 27186 6466 27198
rect 6414 27122 6466 27134
rect 8878 27186 8930 27198
rect 8878 27122 8930 27134
rect 9214 27186 9266 27198
rect 9214 27122 9266 27134
rect 10558 27186 10610 27198
rect 14142 27186 14194 27198
rect 12562 27134 12574 27186
rect 12626 27134 12638 27186
rect 10558 27122 10610 27134
rect 14142 27122 14194 27134
rect 15262 27186 15314 27198
rect 15262 27122 15314 27134
rect 17166 27186 17218 27198
rect 17166 27122 17218 27134
rect 18062 27186 18114 27198
rect 18062 27122 18114 27134
rect 18510 27186 18562 27198
rect 18510 27122 18562 27134
rect 19406 27186 19458 27198
rect 19406 27122 19458 27134
rect 20190 27186 20242 27198
rect 20190 27122 20242 27134
rect 23774 27186 23826 27198
rect 23774 27122 23826 27134
rect 27134 27186 27186 27198
rect 27134 27122 27186 27134
rect 4286 27074 4338 27086
rect 3938 27022 3950 27074
rect 4002 27022 4014 27074
rect 4286 27010 4338 27022
rect 5854 27074 5906 27086
rect 5854 27010 5906 27022
rect 9102 27074 9154 27086
rect 9102 27010 9154 27022
rect 9774 27074 9826 27086
rect 9774 27010 9826 27022
rect 14478 27074 14530 27086
rect 14478 27010 14530 27022
rect 14702 27074 14754 27086
rect 14702 27010 14754 27022
rect 15150 27074 15202 27086
rect 15150 27010 15202 27022
rect 15710 27074 15762 27086
rect 15710 27010 15762 27022
rect 16046 27074 16098 27086
rect 16046 27010 16098 27022
rect 18622 27074 18674 27086
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 24434 27022 24446 27074
rect 24498 27022 24510 27074
rect 25218 27022 25230 27074
rect 25282 27022 25294 27074
rect 26002 27022 26014 27074
rect 26066 27022 26078 27074
rect 18622 27010 18674 27022
rect 3502 26962 3554 26974
rect 3502 26898 3554 26910
rect 8094 26962 8146 26974
rect 8094 26898 8146 26910
rect 10110 26962 10162 26974
rect 10110 26898 10162 26910
rect 12126 26962 12178 26974
rect 12126 26898 12178 26910
rect 13582 26962 13634 26974
rect 13582 26898 13634 26910
rect 15374 26962 15426 26974
rect 15374 26898 15426 26910
rect 15822 26962 15874 26974
rect 15822 26898 15874 26910
rect 17614 26962 17666 26974
rect 17614 26898 17666 26910
rect 18398 26962 18450 26974
rect 18398 26898 18450 26910
rect 18846 26962 18898 26974
rect 25778 26910 25790 26962
rect 25842 26910 25854 26962
rect 18846 26898 18898 26910
rect 3726 26850 3778 26862
rect 3726 26786 3778 26798
rect 9326 26850 9378 26862
rect 9326 26786 9378 26798
rect 16606 26850 16658 26862
rect 16606 26786 16658 26798
rect 21982 26850 22034 26862
rect 21982 26786 22034 26798
rect 26574 26850 26626 26862
rect 26574 26786 26626 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 9662 26514 9714 26526
rect 9662 26450 9714 26462
rect 9774 26514 9826 26526
rect 9774 26450 9826 26462
rect 10558 26514 10610 26526
rect 10558 26450 10610 26462
rect 11006 26514 11058 26526
rect 11006 26450 11058 26462
rect 12798 26514 12850 26526
rect 12798 26450 12850 26462
rect 13246 26514 13298 26526
rect 13246 26450 13298 26462
rect 13694 26514 13746 26526
rect 13694 26450 13746 26462
rect 14142 26514 14194 26526
rect 14142 26450 14194 26462
rect 14702 26514 14754 26526
rect 14702 26450 14754 26462
rect 15598 26514 15650 26526
rect 15598 26450 15650 26462
rect 17726 26514 17778 26526
rect 17726 26450 17778 26462
rect 19518 26514 19570 26526
rect 19518 26450 19570 26462
rect 20414 26514 20466 26526
rect 20414 26450 20466 26462
rect 21758 26514 21810 26526
rect 21758 26450 21810 26462
rect 26014 26514 26066 26526
rect 26014 26450 26066 26462
rect 26574 26514 26626 26526
rect 26574 26450 26626 26462
rect 7646 26402 7698 26414
rect 7646 26338 7698 26350
rect 7870 26402 7922 26414
rect 7870 26338 7922 26350
rect 15038 26402 15090 26414
rect 15038 26338 15090 26350
rect 15710 26402 15762 26414
rect 15710 26338 15762 26350
rect 17614 26402 17666 26414
rect 17614 26338 17666 26350
rect 20862 26402 20914 26414
rect 20862 26338 20914 26350
rect 5518 26290 5570 26302
rect 7310 26290 7362 26302
rect 5954 26238 5966 26290
rect 6018 26238 6030 26290
rect 5518 26226 5570 26238
rect 7310 26226 7362 26238
rect 8206 26290 8258 26302
rect 8206 26226 8258 26238
rect 9550 26290 9602 26302
rect 11342 26290 11394 26302
rect 10098 26238 10110 26290
rect 10162 26238 10174 26290
rect 9550 26226 9602 26238
rect 11342 26226 11394 26238
rect 11902 26290 11954 26302
rect 11902 26226 11954 26238
rect 12238 26290 12290 26302
rect 12238 26226 12290 26238
rect 15486 26290 15538 26302
rect 15486 26226 15538 26238
rect 15822 26290 15874 26302
rect 17838 26290 17890 26302
rect 16034 26238 16046 26290
rect 16098 26238 16110 26290
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 15822 26226 15874 26238
rect 17838 26226 17890 26238
rect 17950 26290 18002 26302
rect 17950 26226 18002 26238
rect 18510 26290 18562 26302
rect 18510 26226 18562 26238
rect 21198 26290 21250 26302
rect 21198 26226 21250 26238
rect 22206 26290 22258 26302
rect 22206 26226 22258 26238
rect 8766 26178 8818 26190
rect 8766 26114 8818 26126
rect 16830 26178 16882 26190
rect 16830 26114 16882 26126
rect 19070 26178 19122 26190
rect 19070 26114 19122 26126
rect 19966 26178 20018 26190
rect 19966 26114 20018 26126
rect 22766 26178 22818 26190
rect 22766 26114 22818 26126
rect 23214 26178 23266 26190
rect 23214 26114 23266 26126
rect 25454 26178 25506 26190
rect 25454 26114 25506 26126
rect 7086 26066 7138 26078
rect 7086 26002 7138 26014
rect 7758 26066 7810 26078
rect 7758 26002 7810 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 8206 25618 8258 25630
rect 7298 25566 7310 25618
rect 7362 25566 7374 25618
rect 8206 25554 8258 25566
rect 8542 25618 8594 25630
rect 8542 25554 8594 25566
rect 14926 25618 14978 25630
rect 27134 25618 27186 25630
rect 29262 25618 29314 25630
rect 16482 25566 16494 25618
rect 16546 25566 16558 25618
rect 17714 25566 17726 25618
rect 17778 25566 17790 25618
rect 19954 25566 19966 25618
rect 20018 25566 20030 25618
rect 28242 25566 28254 25618
rect 28306 25566 28318 25618
rect 14926 25554 14978 25566
rect 27134 25554 27186 25566
rect 29262 25554 29314 25566
rect 9438 25506 9490 25518
rect 7634 25454 7646 25506
rect 7698 25454 7710 25506
rect 8978 25454 8990 25506
rect 9042 25454 9054 25506
rect 9438 25442 9490 25454
rect 9662 25506 9714 25518
rect 9662 25442 9714 25454
rect 10222 25506 10274 25518
rect 10222 25442 10274 25454
rect 10446 25506 10498 25518
rect 11790 25506 11842 25518
rect 10994 25454 11006 25506
rect 11058 25454 11070 25506
rect 10446 25442 10498 25454
rect 11790 25442 11842 25454
rect 11902 25506 11954 25518
rect 12910 25506 12962 25518
rect 12338 25454 12350 25506
rect 12402 25454 12414 25506
rect 14242 25454 14254 25506
rect 14306 25454 14318 25506
rect 15250 25454 15262 25506
rect 15314 25454 15326 25506
rect 16034 25454 16046 25506
rect 16098 25454 16110 25506
rect 17378 25454 17390 25506
rect 17442 25454 17454 25506
rect 18162 25454 18174 25506
rect 18226 25454 18238 25506
rect 18834 25454 18846 25506
rect 18898 25454 18910 25506
rect 19282 25454 19294 25506
rect 19346 25454 19358 25506
rect 20066 25454 20078 25506
rect 20130 25454 20142 25506
rect 21746 25454 21758 25506
rect 21810 25454 21822 25506
rect 23650 25454 23662 25506
rect 23714 25454 23726 25506
rect 25218 25454 25230 25506
rect 25282 25454 25294 25506
rect 25554 25454 25566 25506
rect 25618 25454 25630 25506
rect 27906 25454 27918 25506
rect 27970 25454 27982 25506
rect 11902 25442 11954 25454
rect 12910 25442 12962 25454
rect 1710 25394 1762 25406
rect 1710 25330 1762 25342
rect 2046 25394 2098 25406
rect 2046 25330 2098 25342
rect 2494 25394 2546 25406
rect 2494 25330 2546 25342
rect 6862 25394 6914 25406
rect 6862 25330 6914 25342
rect 9550 25394 9602 25406
rect 9550 25330 9602 25342
rect 10782 25394 10834 25406
rect 10782 25330 10834 25342
rect 12574 25394 12626 25406
rect 14018 25342 14030 25394
rect 14082 25342 14094 25394
rect 16370 25342 16382 25394
rect 16434 25342 16446 25394
rect 17602 25342 17614 25394
rect 17666 25342 17678 25394
rect 20402 25342 20414 25394
rect 20466 25342 20478 25394
rect 22530 25342 22542 25394
rect 22594 25342 22606 25394
rect 23538 25342 23550 25394
rect 23602 25342 23614 25394
rect 12574 25330 12626 25342
rect 9886 25282 9938 25294
rect 12014 25282 12066 25294
rect 11330 25230 11342 25282
rect 11394 25230 11406 25282
rect 9886 25218 9938 25230
rect 12014 25218 12066 25230
rect 12798 25282 12850 25294
rect 12798 25218 12850 25230
rect 13694 25282 13746 25294
rect 21534 25282 21586 25294
rect 15250 25230 15262 25282
rect 15314 25230 15326 25282
rect 18610 25230 18622 25282
rect 18674 25230 18686 25282
rect 21858 25230 21870 25282
rect 21922 25230 21934 25282
rect 13694 25218 13746 25230
rect 21534 25218 21586 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 11230 24946 11282 24958
rect 11230 24882 11282 24894
rect 11678 24946 11730 24958
rect 17614 24946 17666 24958
rect 16706 24894 16718 24946
rect 16770 24894 16782 24946
rect 22978 24894 22990 24946
rect 23042 24894 23054 24946
rect 11678 24882 11730 24894
rect 17614 24882 17666 24894
rect 16034 24782 16046 24834
rect 16098 24782 16110 24834
rect 19282 24782 19294 24834
rect 19346 24782 19358 24834
rect 20402 24782 20414 24834
rect 20466 24782 20478 24834
rect 22418 24782 22430 24834
rect 22482 24782 22494 24834
rect 24210 24782 24222 24834
rect 24274 24782 24286 24834
rect 25790 24722 25842 24734
rect 13010 24670 13022 24722
rect 13074 24670 13086 24722
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 13570 24670 13582 24722
rect 13634 24670 13646 24722
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 16482 24670 16494 24722
rect 16546 24670 16558 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 21074 24670 21086 24722
rect 21138 24670 21150 24722
rect 21970 24670 21982 24722
rect 22034 24670 22046 24722
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 25790 24658 25842 24670
rect 26238 24610 26290 24622
rect 19170 24558 19182 24610
rect 19234 24558 19246 24610
rect 25330 24558 25342 24610
rect 25394 24558 25406 24610
rect 26238 24546 26290 24558
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 20738 24110 20750 24162
rect 20802 24110 20814 24162
rect 11678 24050 11730 24062
rect 16158 24050 16210 24062
rect 21534 24050 21586 24062
rect 24222 24050 24274 24062
rect 12450 23998 12462 24050
rect 12514 23998 12526 24050
rect 14018 23998 14030 24050
rect 14082 23998 14094 24050
rect 15138 23998 15150 24050
rect 15202 23998 15214 24050
rect 19730 23998 19742 24050
rect 19794 23998 19806 24050
rect 23426 23998 23438 24050
rect 23490 23998 23502 24050
rect 11678 23986 11730 23998
rect 16158 23986 16210 23998
rect 21534 23986 21586 23998
rect 24222 23986 24274 23998
rect 25230 24050 25282 24062
rect 25230 23986 25282 23998
rect 25790 24050 25842 24062
rect 25790 23986 25842 23998
rect 12910 23938 12962 23950
rect 15598 23938 15650 23950
rect 20190 23938 20242 23950
rect 14690 23886 14702 23938
rect 14754 23886 14766 23938
rect 16370 23886 16382 23938
rect 16434 23886 16446 23938
rect 17938 23886 17950 23938
rect 18002 23886 18014 23938
rect 19954 23886 19966 23938
rect 20018 23886 20030 23938
rect 12910 23874 12962 23886
rect 15598 23874 15650 23886
rect 20190 23874 20242 23886
rect 20302 23938 20354 23950
rect 24782 23938 24834 23950
rect 21970 23886 21982 23938
rect 22034 23886 22046 23938
rect 22306 23886 22318 23938
rect 22370 23886 22382 23938
rect 23762 23886 23774 23938
rect 23826 23886 23838 23938
rect 20302 23874 20354 23886
rect 24782 23874 24834 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 2046 23826 2098 23838
rect 16930 23774 16942 23826
rect 16994 23774 17006 23826
rect 18162 23774 18174 23826
rect 18226 23774 18238 23826
rect 21298 23774 21310 23826
rect 21362 23774 21374 23826
rect 2046 23762 2098 23774
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 15150 23378 15202 23390
rect 15150 23314 15202 23326
rect 15598 23378 15650 23390
rect 15598 23314 15650 23326
rect 15934 23378 15986 23390
rect 15934 23314 15986 23326
rect 16158 23378 16210 23390
rect 16158 23314 16210 23326
rect 16606 23378 16658 23390
rect 16606 23314 16658 23326
rect 19070 23378 19122 23390
rect 19070 23314 19122 23326
rect 21086 23378 21138 23390
rect 21086 23314 21138 23326
rect 21646 23378 21698 23390
rect 21646 23314 21698 23326
rect 22990 23378 23042 23390
rect 22990 23314 23042 23326
rect 25454 23378 25506 23390
rect 25454 23314 25506 23326
rect 15822 23266 15874 23278
rect 15822 23202 15874 23214
rect 19182 23266 19234 23278
rect 22206 23266 22258 23278
rect 21298 23214 21310 23266
rect 21362 23214 21374 23266
rect 19182 23202 19234 23214
rect 22206 23202 22258 23214
rect 17614 23042 17666 23054
rect 17614 22978 17666 22990
rect 19070 22930 19122 22942
rect 19070 22866 19122 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 1710 22258 1762 22270
rect 1710 22194 1762 22206
rect 2046 22258 2098 22270
rect 2046 22194 2098 22206
rect 2494 22146 2546 22158
rect 2494 22082 2546 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 2034 20638 2046 20690
rect 2098 20638 2110 20690
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 2494 20578 2546 20590
rect 2494 20514 2546 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 2046 18674 2098 18686
rect 2046 18610 2098 18622
rect 1710 18450 1762 18462
rect 1710 18386 1762 18398
rect 2494 18338 2546 18350
rect 2494 18274 2546 18286
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 2034 17054 2046 17106
rect 2098 17054 2110 17106
rect 1710 16882 1762 16894
rect 1710 16818 1762 16830
rect 2494 16882 2546 16894
rect 2494 16818 2546 16830
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 2046 15538 2098 15550
rect 2046 15474 2098 15486
rect 1710 15314 1762 15326
rect 1710 15250 1762 15262
rect 2494 15202 2546 15214
rect 2494 15138 2546 15150
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 2046 12850 2098 12862
rect 2046 12786 2098 12798
rect 2494 12850 2546 12862
rect 2494 12786 2546 12798
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 1710 11282 1762 11294
rect 1710 11218 1762 11230
rect 2046 11282 2098 11294
rect 2046 11218 2098 11230
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 2494 9602 2546 9614
rect 2494 9538 2546 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2046 8146 2098 8158
rect 2046 8082 2098 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 1710 5906 1762 5918
rect 1710 5842 1762 5854
rect 2146 5742 2158 5794
rect 2210 5742 2222 5794
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 1822 5234 1874 5246
rect 1822 5170 1874 5182
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 2046 4562 2098 4574
rect 2046 4498 2098 4510
rect 1710 4338 1762 4350
rect 1710 4274 1762 4286
rect 2494 4226 2546 4238
rect 2494 4162 2546 4174
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 2270 3666 2322 3678
rect 2270 3602 2322 3614
rect 1710 3442 1762 3454
rect 1710 3378 1762 3390
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 38782 56590 38834 56642
rect 39342 56590 39394 56642
rect 40126 56590 40178 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 5070 56254 5122 56306
rect 7422 56254 7474 56306
rect 7646 56254 7698 56306
rect 9662 56254 9714 56306
rect 9886 56254 9938 56306
rect 11902 56254 11954 56306
rect 12126 56254 12178 56306
rect 14142 56254 14194 56306
rect 16494 56254 16546 56306
rect 16942 56254 16994 56306
rect 18622 56254 18674 56306
rect 18846 56254 18898 56306
rect 20302 56254 20354 56306
rect 23102 56254 23154 56306
rect 25342 56254 25394 56306
rect 29822 56254 29874 56306
rect 31726 56254 31778 56306
rect 34302 56254 34354 56306
rect 36542 56254 36594 56306
rect 39342 56254 39394 56306
rect 41470 56254 41522 56306
rect 44606 56254 44658 56306
rect 48974 56254 49026 56306
rect 52222 56254 52274 56306
rect 56030 56254 56082 56306
rect 2046 56142 2098 56194
rect 2382 56142 2434 56194
rect 5518 56142 5570 56194
rect 5854 56142 5906 56194
rect 7982 56142 8034 56194
rect 10222 56142 10274 56194
rect 12462 56142 12514 56194
rect 14366 56142 14418 56194
rect 17278 56142 17330 56194
rect 19182 56142 19234 56194
rect 21086 56142 21138 56194
rect 21422 56142 21474 56194
rect 23326 56142 23378 56194
rect 25566 56142 25618 56194
rect 28366 56142 28418 56194
rect 30046 56142 30098 56194
rect 32286 56142 32338 56194
rect 32622 56142 32674 56194
rect 34526 56142 34578 56194
rect 34862 56142 34914 56194
rect 36766 56142 36818 56194
rect 37102 56142 37154 56194
rect 39790 56142 39842 56194
rect 40126 56142 40178 56194
rect 1710 56030 1762 56082
rect 2606 56030 2658 56082
rect 14590 56030 14642 56082
rect 23550 56030 23602 56082
rect 25790 56030 25842 56082
rect 28590 56030 28642 56082
rect 30270 56030 30322 56082
rect 40462 56030 40514 56082
rect 43710 56030 43762 56082
rect 47742 56030 47794 56082
rect 47966 56030 48018 56082
rect 51214 56030 51266 56082
rect 54574 56030 54626 56082
rect 55022 56030 55074 56082
rect 3166 55918 3218 55970
rect 27918 55918 27970 55970
rect 38894 55918 38946 55970
rect 27582 55806 27634 55858
rect 27918 55806 27970 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 2158 55358 2210 55410
rect 16382 55358 16434 55410
rect 20526 55358 20578 55410
rect 32062 55358 32114 55410
rect 36430 55358 36482 55410
rect 39118 55358 39170 55410
rect 43150 55358 43202 55410
rect 46734 55358 46786 55410
rect 53678 55358 53730 55410
rect 56702 55358 56754 55410
rect 13582 55246 13634 55298
rect 16830 55246 16882 55298
rect 17726 55246 17778 55298
rect 21422 55246 21474 55298
rect 22990 55246 23042 55298
rect 25454 55246 25506 55298
rect 27694 55246 27746 55298
rect 29262 55246 29314 55298
rect 32622 55246 32674 55298
rect 33630 55246 33682 55298
rect 37102 55246 37154 55298
rect 38334 55246 38386 55298
rect 40238 55246 40290 55298
rect 45726 55246 45778 55298
rect 52670 55246 52722 55298
rect 55582 55246 55634 55298
rect 11790 55134 11842 55186
rect 14254 55134 14306 55186
rect 18398 55134 18450 55186
rect 29934 55134 29986 55186
rect 34302 55134 34354 55186
rect 37326 55134 37378 55186
rect 41022 55134 41074 55186
rect 11902 55022 11954 55074
rect 22878 55022 22930 55074
rect 25342 55022 25394 55074
rect 27582 55022 27634 55074
rect 32622 55022 32674 55074
rect 33182 55022 33234 55074
rect 37774 55022 37826 55074
rect 38110 55022 38162 55074
rect 39006 55022 39058 55074
rect 39902 55022 39954 55074
rect 43598 55022 43650 55074
rect 45390 55022 45442 55074
rect 50878 55022 50930 55074
rect 52110 55022 52162 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 14702 54686 14754 54738
rect 15822 54686 15874 54738
rect 17614 54686 17666 54738
rect 18510 54686 18562 54738
rect 29486 54686 29538 54738
rect 29934 54686 29986 54738
rect 32510 54686 32562 54738
rect 33966 54686 34018 54738
rect 41022 54686 41074 54738
rect 2046 54574 2098 54626
rect 12798 54574 12850 54626
rect 13134 54574 13186 54626
rect 15150 54574 15202 54626
rect 29150 54574 29202 54626
rect 31838 54574 31890 54626
rect 33406 54574 33458 54626
rect 36206 54574 36258 54626
rect 38894 54574 38946 54626
rect 39566 54574 39618 54626
rect 40910 54574 40962 54626
rect 1710 54462 1762 54514
rect 12462 54462 12514 54514
rect 13694 54462 13746 54514
rect 14590 54462 14642 54514
rect 14926 54462 14978 54514
rect 15710 54462 15762 54514
rect 15934 54462 15986 54514
rect 16382 54462 16434 54514
rect 17278 54462 17330 54514
rect 17614 54462 17666 54514
rect 17838 54462 17890 54514
rect 18286 54462 18338 54514
rect 18398 54462 18450 54514
rect 18846 54462 18898 54514
rect 20974 54462 21026 54514
rect 25230 54462 25282 54514
rect 28814 54462 28866 54514
rect 29822 54462 29874 54514
rect 30046 54462 30098 54514
rect 30606 54462 30658 54514
rect 33182 54462 33234 54514
rect 33966 54462 34018 54514
rect 34862 54462 34914 54514
rect 38222 54462 38274 54514
rect 38558 54462 38610 54514
rect 39230 54462 39282 54514
rect 41134 54462 41186 54514
rect 41358 54462 41410 54514
rect 41470 54462 41522 54514
rect 2494 54350 2546 54402
rect 13806 54350 13858 54402
rect 21758 54350 21810 54402
rect 23886 54350 23938 54402
rect 26014 54350 26066 54402
rect 28142 54350 28194 54402
rect 31726 54350 31778 54402
rect 34750 54350 34802 54402
rect 36094 54350 36146 54402
rect 36878 54350 36930 54402
rect 40350 54350 40402 54402
rect 55246 54350 55298 54402
rect 30382 54238 30434 54290
rect 32062 54238 32114 54290
rect 33630 54238 33682 54290
rect 36430 54238 36482 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 40910 53902 40962 53954
rect 41246 53902 41298 53954
rect 23662 53790 23714 53842
rect 26350 53790 26402 53842
rect 29262 53790 29314 53842
rect 37662 53790 37714 53842
rect 38894 53790 38946 53842
rect 42030 53790 42082 53842
rect 16382 53678 16434 53730
rect 18174 53678 18226 53730
rect 21982 53678 22034 53730
rect 22430 53678 22482 53730
rect 22654 53678 22706 53730
rect 22878 53678 22930 53730
rect 24446 53678 24498 53730
rect 25118 53678 25170 53730
rect 33070 53678 33122 53730
rect 38222 53678 38274 53730
rect 41246 53678 41298 53730
rect 16606 53566 16658 53618
rect 22318 53566 22370 53618
rect 24894 53566 24946 53618
rect 32622 53566 32674 53618
rect 33294 53566 33346 53618
rect 42366 53566 42418 53618
rect 10446 53454 10498 53506
rect 11566 53454 11618 53506
rect 15374 53454 15426 53506
rect 15934 53454 15986 53506
rect 23550 53454 23602 53506
rect 23774 53454 23826 53506
rect 23998 53454 24050 53506
rect 24782 53454 24834 53506
rect 25566 53454 25618 53506
rect 26238 53454 26290 53506
rect 26462 53454 26514 53506
rect 26686 53454 26738 53506
rect 37998 53454 38050 53506
rect 42142 53454 42194 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 12798 53118 12850 53170
rect 23438 53118 23490 53170
rect 29150 53118 29202 53170
rect 31950 53118 32002 53170
rect 33854 53118 33906 53170
rect 41358 53118 41410 53170
rect 2046 53006 2098 53058
rect 7982 53006 8034 53058
rect 9886 53006 9938 53058
rect 10670 53006 10722 53058
rect 12014 53006 12066 53058
rect 12350 53006 12402 53058
rect 22766 53006 22818 53058
rect 26686 53006 26738 53058
rect 29598 53006 29650 53058
rect 29934 53006 29986 53058
rect 30158 53006 30210 53058
rect 32174 53006 32226 53058
rect 33070 53006 33122 53058
rect 36430 53006 36482 53058
rect 36542 53006 36594 53058
rect 40910 53006 40962 53058
rect 42814 53006 42866 53058
rect 1710 52894 1762 52946
rect 8766 52894 8818 52946
rect 10222 52894 10274 52946
rect 10558 52894 10610 52946
rect 10894 52894 10946 52946
rect 11342 52894 11394 52946
rect 17950 52894 18002 52946
rect 18398 52894 18450 52946
rect 18510 52894 18562 52946
rect 22318 52894 22370 52946
rect 22990 52894 23042 52946
rect 25454 52894 25506 52946
rect 25902 52894 25954 52946
rect 26126 52894 26178 52946
rect 27022 52894 27074 52946
rect 30382 52894 30434 52946
rect 30718 52894 30770 52946
rect 33294 52894 33346 52946
rect 33854 52894 33906 52946
rect 36766 52894 36818 52946
rect 41134 52894 41186 52946
rect 41694 52894 41746 52946
rect 42030 52894 42082 52946
rect 2494 52782 2546 52834
rect 5854 52782 5906 52834
rect 15374 52782 15426 52834
rect 18174 52782 18226 52834
rect 19070 52782 19122 52834
rect 22542 52782 22594 52834
rect 26014 52782 26066 52834
rect 27470 52782 27522 52834
rect 30046 52782 30098 52834
rect 31838 52782 31890 52834
rect 36206 52782 36258 52834
rect 40350 52782 40402 52834
rect 44942 52782 44994 52834
rect 2270 52670 2322 52722
rect 2606 52670 2658 52722
rect 11006 52670 11058 52722
rect 25118 52670 25170 52722
rect 25342 52670 25394 52722
rect 29486 52670 29538 52722
rect 33630 52670 33682 52722
rect 37214 52670 37266 52722
rect 41470 52670 41522 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 10446 52334 10498 52386
rect 11678 52334 11730 52386
rect 12798 52222 12850 52274
rect 15598 52222 15650 52274
rect 17838 52222 17890 52274
rect 19966 52222 20018 52274
rect 22094 52222 22146 52274
rect 30158 52222 30210 52274
rect 32286 52222 32338 52274
rect 32734 52222 32786 52274
rect 34078 52222 34130 52274
rect 36206 52222 36258 52274
rect 36990 52222 37042 52274
rect 37102 52222 37154 52274
rect 38670 52222 38722 52274
rect 41246 52222 41298 52274
rect 42590 52222 42642 52274
rect 8990 52110 9042 52162
rect 9998 52110 10050 52162
rect 10334 52110 10386 52162
rect 10782 52110 10834 52162
rect 11118 52110 11170 52162
rect 11342 52110 11394 52162
rect 11902 52110 11954 52162
rect 12350 52110 12402 52162
rect 14590 52110 14642 52162
rect 14814 52110 14866 52162
rect 15150 52110 15202 52162
rect 15710 52110 15762 52162
rect 16046 52110 16098 52162
rect 20750 52110 20802 52162
rect 27022 52110 27074 52162
rect 27470 52110 27522 52162
rect 29374 52110 29426 52162
rect 33406 52110 33458 52162
rect 37326 52110 37378 52162
rect 38222 52110 38274 52162
rect 40238 52110 40290 52162
rect 42478 52110 42530 52162
rect 42926 52110 42978 52162
rect 39118 51998 39170 52050
rect 42142 51998 42194 52050
rect 10110 51886 10162 51938
rect 11902 51886 11954 51938
rect 14702 51886 14754 51938
rect 15486 51886 15538 51938
rect 41694 51886 41746 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 12014 51550 12066 51602
rect 16494 51550 16546 51602
rect 23102 51550 23154 51602
rect 38894 51550 38946 51602
rect 40126 51550 40178 51602
rect 42254 51550 42306 51602
rect 2046 51438 2098 51490
rect 10670 51438 10722 51490
rect 10894 51438 10946 51490
rect 13918 51438 13970 51490
rect 18734 51438 18786 51490
rect 39678 51438 39730 51490
rect 40350 51438 40402 51490
rect 41022 51438 41074 51490
rect 41246 51438 41298 51490
rect 1822 51326 1874 51378
rect 4398 51326 4450 51378
rect 7646 51326 7698 51378
rect 11118 51326 11170 51378
rect 11230 51326 11282 51378
rect 13134 51326 13186 51378
rect 16830 51326 16882 51378
rect 22654 51326 22706 51378
rect 25342 51326 25394 51378
rect 39118 51326 39170 51378
rect 39454 51326 39506 51378
rect 41470 51326 41522 51378
rect 41806 51326 41858 51378
rect 2494 51214 2546 51266
rect 5070 51214 5122 51266
rect 7198 51214 7250 51266
rect 10782 51214 10834 51266
rect 16046 51214 16098 51266
rect 26126 51214 26178 51266
rect 28254 51214 28306 51266
rect 36430 51214 36482 51266
rect 38558 51214 38610 51266
rect 41134 51214 41186 51266
rect 42142 51214 42194 51266
rect 39230 51102 39282 51154
rect 40014 51102 40066 51154
rect 42478 51102 42530 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 7310 50766 7362 50818
rect 1710 50654 1762 50706
rect 3838 50654 3890 50706
rect 5070 50654 5122 50706
rect 7086 50654 7138 50706
rect 15934 50654 15986 50706
rect 16494 50654 16546 50706
rect 18286 50654 18338 50706
rect 22094 50654 22146 50706
rect 24222 50654 24274 50706
rect 26462 50654 26514 50706
rect 27358 50654 27410 50706
rect 34638 50654 34690 50706
rect 37998 50654 38050 50706
rect 40126 50654 40178 50706
rect 44158 50654 44210 50706
rect 4622 50542 4674 50594
rect 17390 50542 17442 50594
rect 18174 50542 18226 50594
rect 18846 50542 18898 50594
rect 21422 50542 21474 50594
rect 25230 50542 25282 50594
rect 26238 50542 26290 50594
rect 26686 50542 26738 50594
rect 26798 50542 26850 50594
rect 30270 50542 30322 50594
rect 35198 50542 35250 50594
rect 36430 50542 36482 50594
rect 37326 50542 37378 50594
rect 40910 50542 40962 50594
rect 41358 50542 41410 50594
rect 17726 50430 17778 50482
rect 18398 50430 18450 50482
rect 24782 50430 24834 50482
rect 25454 50430 25506 50482
rect 42030 50430 42082 50482
rect 7646 50318 7698 50370
rect 11902 50318 11954 50370
rect 12574 50318 12626 50370
rect 16046 50318 16098 50370
rect 24558 50318 24610 50370
rect 24670 50318 24722 50370
rect 25790 50318 25842 50370
rect 30606 50318 30658 50370
rect 32398 50318 32450 50370
rect 34974 50318 35026 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 5070 49982 5122 50034
rect 11342 49982 11394 50034
rect 12014 49982 12066 50034
rect 15262 49982 15314 50034
rect 22430 49982 22482 50034
rect 33182 49982 33234 50034
rect 3838 49870 3890 49922
rect 7198 49870 7250 49922
rect 7534 49870 7586 49922
rect 13134 49870 13186 49922
rect 25230 49870 25282 49922
rect 27582 49870 27634 49922
rect 4622 49758 4674 49810
rect 6526 49758 6578 49810
rect 8878 49758 8930 49810
rect 10446 49758 10498 49810
rect 11566 49758 11618 49810
rect 12238 49758 12290 49810
rect 12910 49758 12962 49810
rect 22094 49758 22146 49810
rect 32174 49758 32226 49810
rect 37326 49758 37378 49810
rect 1710 49646 1762 49698
rect 6414 49646 6466 49698
rect 6974 49646 7026 49698
rect 7982 49646 8034 49698
rect 8542 49646 8594 49698
rect 10110 49646 10162 49698
rect 14926 49646 14978 49698
rect 21758 49646 21810 49698
rect 25790 49646 25842 49698
rect 29262 49646 29314 49698
rect 31390 49646 31442 49698
rect 34414 49646 34466 49698
rect 36542 49646 36594 49698
rect 37774 49646 37826 49698
rect 11230 49534 11282 49586
rect 11902 49534 11954 49586
rect 25342 49534 25394 49586
rect 27694 49534 27746 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 35870 49198 35922 49250
rect 36542 49198 36594 49250
rect 6638 49086 6690 49138
rect 10222 49086 10274 49138
rect 11342 49086 11394 49138
rect 11902 49086 11954 49138
rect 12462 49086 12514 49138
rect 14366 49086 14418 49138
rect 15934 49086 15986 49138
rect 19182 49086 19234 49138
rect 19966 49086 20018 49138
rect 24558 49086 24610 49138
rect 29598 49086 29650 49138
rect 35534 49086 35586 49138
rect 38446 49086 38498 49138
rect 7086 48974 7138 49026
rect 11454 48974 11506 49026
rect 13918 48974 13970 49026
rect 14142 48974 14194 49026
rect 15150 48974 15202 49026
rect 15374 48974 15426 49026
rect 16494 48974 16546 49026
rect 17502 48974 17554 49026
rect 18062 48974 18114 49026
rect 19070 48974 19122 49026
rect 19406 48974 19458 49026
rect 20526 48974 20578 49026
rect 21870 48974 21922 49026
rect 22094 48974 22146 49026
rect 22206 48974 22258 49026
rect 24670 48974 24722 49026
rect 25678 48974 25730 49026
rect 27134 48974 27186 49026
rect 27918 48974 27970 49026
rect 32510 48974 32562 49026
rect 32846 48974 32898 49026
rect 34190 48974 34242 49026
rect 34302 48974 34354 49026
rect 35086 48974 35138 49026
rect 35422 48974 35474 49026
rect 1710 48862 1762 48914
rect 11118 48862 11170 48914
rect 16382 48862 16434 48914
rect 17614 48862 17666 48914
rect 17838 48862 17890 48914
rect 19630 48862 19682 48914
rect 19854 48862 19906 48914
rect 20414 48862 20466 48914
rect 22542 48862 22594 48914
rect 22878 48862 22930 48914
rect 22990 48862 23042 48914
rect 25454 48862 25506 48914
rect 27358 48862 27410 48914
rect 31726 48862 31778 48914
rect 33070 48862 33122 48914
rect 35646 48862 35698 48914
rect 2046 48750 2098 48802
rect 2494 48750 2546 48802
rect 9662 48750 9714 48802
rect 13470 48750 13522 48802
rect 14814 48750 14866 48802
rect 16158 48750 16210 48802
rect 18398 48750 18450 48802
rect 18846 48750 18898 48802
rect 20190 48750 20242 48802
rect 22430 48750 22482 48802
rect 23214 48750 23266 48802
rect 32958 48750 33010 48802
rect 33294 48750 33346 48802
rect 33854 48750 33906 48802
rect 34414 48750 34466 48802
rect 34638 48750 34690 48802
rect 36094 48750 36146 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 3502 48414 3554 48466
rect 16270 48414 16322 48466
rect 16718 48414 16770 48466
rect 17950 48414 18002 48466
rect 19966 48414 20018 48466
rect 30494 48414 30546 48466
rect 31390 48414 31442 48466
rect 38782 48414 38834 48466
rect 7086 48302 7138 48354
rect 10558 48302 10610 48354
rect 12126 48302 12178 48354
rect 15710 48302 15762 48354
rect 17502 48302 17554 48354
rect 19182 48302 19234 48354
rect 19854 48302 19906 48354
rect 21534 48302 21586 48354
rect 21870 48302 21922 48354
rect 22878 48302 22930 48354
rect 23438 48302 23490 48354
rect 23886 48302 23938 48354
rect 23998 48302 24050 48354
rect 26462 48302 26514 48354
rect 27358 48302 27410 48354
rect 29822 48302 29874 48354
rect 30830 48302 30882 48354
rect 31726 48302 31778 48354
rect 39118 48302 39170 48354
rect 6638 48190 6690 48242
rect 7198 48190 7250 48242
rect 9662 48190 9714 48242
rect 10670 48190 10722 48242
rect 11342 48190 11394 48242
rect 11790 48190 11842 48242
rect 13582 48190 13634 48242
rect 13806 48190 13858 48242
rect 14478 48190 14530 48242
rect 15374 48190 15426 48242
rect 18062 48190 18114 48242
rect 20078 48190 20130 48242
rect 22766 48190 22818 48242
rect 23102 48190 23154 48242
rect 23326 48190 23378 48242
rect 23662 48190 23714 48242
rect 24558 48190 24610 48242
rect 26574 48190 26626 48242
rect 27134 48190 27186 48242
rect 28702 48190 28754 48242
rect 29038 48190 29090 48242
rect 31166 48190 31218 48242
rect 31502 48190 31554 48242
rect 33630 48190 33682 48242
rect 4062 48078 4114 48130
rect 6078 48078 6130 48130
rect 10222 48078 10274 48130
rect 13358 48078 13410 48130
rect 15262 48078 15314 48130
rect 18286 48078 18338 48130
rect 20526 48078 20578 48130
rect 22430 48078 22482 48130
rect 32174 48078 32226 48130
rect 38222 48078 38274 48130
rect 39678 48078 39730 48130
rect 7086 47966 7138 48018
rect 14030 47966 14082 48018
rect 17390 47966 17442 48018
rect 22206 47966 22258 48018
rect 22542 47966 22594 48018
rect 23998 47966 24050 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 3278 47630 3330 47682
rect 18622 47630 18674 47682
rect 3054 47518 3106 47570
rect 8766 47518 8818 47570
rect 28254 47518 28306 47570
rect 32062 47518 32114 47570
rect 33070 47518 33122 47570
rect 35646 47518 35698 47570
rect 40014 47518 40066 47570
rect 2158 47406 2210 47458
rect 2718 47406 2770 47458
rect 3950 47406 4002 47458
rect 6638 47406 6690 47458
rect 7870 47406 7922 47458
rect 8318 47406 8370 47458
rect 10670 47406 10722 47458
rect 11118 47406 11170 47458
rect 14926 47406 14978 47458
rect 15262 47406 15314 47458
rect 17166 47406 17218 47458
rect 18286 47406 18338 47458
rect 18398 47406 18450 47458
rect 19182 47406 19234 47458
rect 20078 47406 20130 47458
rect 20302 47406 20354 47458
rect 25566 47406 25618 47458
rect 27470 47406 27522 47458
rect 29598 47406 29650 47458
rect 30942 47406 30994 47458
rect 31278 47406 31330 47458
rect 33742 47406 33794 47458
rect 34862 47406 34914 47458
rect 35198 47406 35250 47458
rect 38110 47406 38162 47458
rect 38558 47406 38610 47458
rect 39006 47406 39058 47458
rect 42814 47406 42866 47458
rect 4510 47294 4562 47346
rect 6190 47294 6242 47346
rect 7310 47294 7362 47346
rect 9214 47294 9266 47346
rect 12798 47294 12850 47346
rect 14030 47294 14082 47346
rect 17278 47294 17330 47346
rect 18734 47294 18786 47346
rect 19406 47294 19458 47346
rect 19854 47294 19906 47346
rect 25790 47294 25842 47346
rect 27806 47294 27858 47346
rect 29150 47294 29202 47346
rect 33406 47294 33458 47346
rect 34638 47294 34690 47346
rect 42142 47294 42194 47346
rect 3614 47182 3666 47234
rect 10110 47182 10162 47234
rect 15038 47182 15090 47234
rect 16494 47182 16546 47234
rect 17502 47182 17554 47234
rect 19294 47182 19346 47234
rect 19742 47182 19794 47234
rect 35086 47182 35138 47234
rect 38782 47182 38834 47234
rect 39454 47182 39506 47234
rect 39566 47182 39618 47234
rect 39678 47182 39730 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 2494 46846 2546 46898
rect 13694 46846 13746 46898
rect 16158 46846 16210 46898
rect 32622 46846 32674 46898
rect 34078 46846 34130 46898
rect 38446 46846 38498 46898
rect 40350 46846 40402 46898
rect 41358 46846 41410 46898
rect 1710 46734 1762 46786
rect 2046 46734 2098 46786
rect 2942 46734 2994 46786
rect 3726 46734 3778 46786
rect 4846 46734 4898 46786
rect 6414 46734 6466 46786
rect 7870 46734 7922 46786
rect 10334 46734 10386 46786
rect 11342 46734 11394 46786
rect 13134 46734 13186 46786
rect 13358 46734 13410 46786
rect 15710 46734 15762 46786
rect 20750 46734 20802 46786
rect 22654 46734 22706 46786
rect 30158 46734 30210 46786
rect 33518 46734 33570 46786
rect 36654 46734 36706 46786
rect 38782 46734 38834 46786
rect 39454 46734 39506 46786
rect 40910 46734 40962 46786
rect 41134 46734 41186 46786
rect 3950 46622 4002 46674
rect 4510 46622 4562 46674
rect 6974 46622 7026 46674
rect 7310 46622 7362 46674
rect 10782 46622 10834 46674
rect 11454 46622 11506 46674
rect 14702 46622 14754 46674
rect 15038 46622 15090 46674
rect 21310 46622 21362 46674
rect 21534 46622 21586 46674
rect 22094 46622 22146 46674
rect 23102 46622 23154 46674
rect 24222 46622 24274 46674
rect 25230 46622 25282 46674
rect 33070 46622 33122 46674
rect 33294 46622 33346 46674
rect 33742 46622 33794 46674
rect 37326 46622 37378 46674
rect 39118 46622 39170 46674
rect 41470 46622 41522 46674
rect 3838 46510 3890 46562
rect 5966 46510 6018 46562
rect 14366 46510 14418 46562
rect 22430 46510 22482 46562
rect 23662 46510 23714 46562
rect 24782 46510 24834 46562
rect 34526 46510 34578 46562
rect 3054 46398 3106 46450
rect 15038 46398 15090 46450
rect 38670 46398 38722 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 33630 46062 33682 46114
rect 9886 45950 9938 46002
rect 14478 45950 14530 46002
rect 17726 45950 17778 46002
rect 22206 45950 22258 46002
rect 26910 45950 26962 46002
rect 32062 45950 32114 46002
rect 32846 45950 32898 46002
rect 33966 45950 34018 46002
rect 34414 45950 34466 46002
rect 41022 45950 41074 46002
rect 3950 45838 4002 45890
rect 6862 45838 6914 45890
rect 7198 45838 7250 45890
rect 7646 45838 7698 45890
rect 8654 45838 8706 45890
rect 10334 45838 10386 45890
rect 12126 45838 12178 45890
rect 13918 45838 13970 45890
rect 15934 45838 15986 45890
rect 16382 45838 16434 45890
rect 16718 45838 16770 45890
rect 17278 45838 17330 45890
rect 19966 45838 20018 45890
rect 20078 45838 20130 45890
rect 21534 45838 21586 45890
rect 21982 45838 22034 45890
rect 24446 45838 24498 45890
rect 24782 45838 24834 45890
rect 26798 45838 26850 45890
rect 29374 45838 29426 45890
rect 30942 45838 30994 45890
rect 31838 45838 31890 45890
rect 32734 45838 32786 45890
rect 32958 45838 33010 45890
rect 34526 45838 34578 45890
rect 41582 45838 41634 45890
rect 41918 45838 41970 45890
rect 1710 45726 1762 45778
rect 4510 45726 4562 45778
rect 6526 45726 6578 45778
rect 9326 45726 9378 45778
rect 10894 45736 10946 45788
rect 16158 45726 16210 45778
rect 21758 45726 21810 45778
rect 22430 45726 22482 45778
rect 23662 45726 23714 45778
rect 24222 45726 24274 45778
rect 24558 45726 24610 45778
rect 24894 45726 24946 45778
rect 27358 45726 27410 45778
rect 29262 45726 29314 45778
rect 33182 45726 33234 45778
rect 34750 45726 34802 45778
rect 41358 45726 41410 45778
rect 2046 45614 2098 45666
rect 2494 45614 2546 45666
rect 6638 45614 6690 45666
rect 8094 45614 8146 45666
rect 10446 45614 10498 45666
rect 16046 45614 16098 45666
rect 19742 45614 19794 45666
rect 20638 45614 20690 45666
rect 22542 45614 22594 45666
rect 33854 45614 33906 45666
rect 34302 45614 34354 45666
rect 38670 45614 38722 45666
rect 41806 45614 41858 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 2606 45278 2658 45330
rect 3166 45278 3218 45330
rect 8206 45278 8258 45330
rect 11230 45278 11282 45330
rect 19742 45278 19794 45330
rect 21422 45278 21474 45330
rect 21646 45278 21698 45330
rect 23326 45278 23378 45330
rect 27582 45278 27634 45330
rect 39230 45278 39282 45330
rect 7982 45166 8034 45218
rect 10670 45166 10722 45218
rect 19070 45166 19122 45218
rect 19406 45166 19458 45218
rect 22318 45166 22370 45218
rect 26238 45166 26290 45218
rect 28702 45166 28754 45218
rect 39006 45166 39058 45218
rect 39342 45166 39394 45218
rect 42366 45166 42418 45218
rect 2494 45054 2546 45106
rect 3054 45054 3106 45106
rect 4174 45054 4226 45106
rect 6862 45054 6914 45106
rect 6974 45054 7026 45106
rect 7758 45054 7810 45106
rect 9774 45054 9826 45106
rect 13694 45054 13746 45106
rect 19966 45054 20018 45106
rect 20750 45054 20802 45106
rect 22094 45054 22146 45106
rect 22206 45054 22258 45106
rect 22766 45054 22818 45106
rect 26126 45054 26178 45106
rect 29822 45054 29874 45106
rect 32510 45054 32562 45106
rect 33406 45054 33458 45106
rect 39566 45054 39618 45106
rect 41582 45054 41634 45106
rect 3726 44942 3778 44994
rect 6750 44942 6802 44994
rect 8206 44942 8258 44994
rect 11454 44942 11506 44994
rect 14254 44942 14306 44994
rect 18622 44942 18674 44994
rect 20302 44942 20354 44994
rect 20526 44942 20578 44994
rect 24670 44942 24722 44994
rect 25342 44942 25394 44994
rect 25790 44942 25842 44994
rect 30382 44942 30434 44994
rect 37102 44942 37154 44994
rect 44494 44942 44546 44994
rect 2606 44830 2658 44882
rect 3166 44830 3218 44882
rect 20974 44830 21026 44882
rect 22990 44830 23042 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 17278 44494 17330 44546
rect 26014 44494 26066 44546
rect 29934 44494 29986 44546
rect 34526 44494 34578 44546
rect 8542 44382 8594 44434
rect 10110 44382 10162 44434
rect 12574 44382 12626 44434
rect 14814 44382 14866 44434
rect 16158 44382 16210 44434
rect 17614 44382 17666 44434
rect 23438 44382 23490 44434
rect 25790 44382 25842 44434
rect 27806 44382 27858 44434
rect 33518 44382 33570 44434
rect 35422 44382 35474 44434
rect 37214 44382 37266 44434
rect 39342 44382 39394 44434
rect 41134 44382 41186 44434
rect 6862 44270 6914 44322
rect 10222 44270 10274 44322
rect 11006 44270 11058 44322
rect 11342 44270 11394 44322
rect 11566 44270 11618 44322
rect 12798 44270 12850 44322
rect 14366 44270 14418 44322
rect 15262 44270 15314 44322
rect 15710 44270 15762 44322
rect 16382 44270 16434 44322
rect 16606 44270 16658 44322
rect 16830 44270 16882 44322
rect 18398 44270 18450 44322
rect 19070 44270 19122 44322
rect 23102 44270 23154 44322
rect 25230 44270 25282 44322
rect 26238 44270 26290 44322
rect 26910 44270 26962 44322
rect 28142 44270 28194 44322
rect 29150 44270 29202 44322
rect 30830 44270 30882 44322
rect 32398 44270 32450 44322
rect 33294 44270 33346 44322
rect 34190 44270 34242 44322
rect 34750 44270 34802 44322
rect 40014 44270 40066 44322
rect 40574 44270 40626 44322
rect 41022 44270 41074 44322
rect 5742 44158 5794 44210
rect 8094 44158 8146 44210
rect 10558 44158 10610 44210
rect 12462 44158 12514 44210
rect 18062 44158 18114 44210
rect 19294 44158 19346 44210
rect 24782 44158 24834 44210
rect 25118 44158 25170 44210
rect 26574 44158 26626 44210
rect 26798 44158 26850 44210
rect 30606 44158 30658 44210
rect 34974 44158 35026 44210
rect 11790 44046 11842 44098
rect 13694 44046 13746 44098
rect 21422 44046 21474 44098
rect 22654 44046 22706 44098
rect 24334 44046 24386 44098
rect 34638 44046 34690 44098
rect 41246 44046 41298 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 17502 43710 17554 43762
rect 22206 43710 22258 43762
rect 29598 43710 29650 43762
rect 39566 43710 39618 43762
rect 41134 43710 41186 43762
rect 3502 43598 3554 43650
rect 5294 43598 5346 43650
rect 6190 43598 6242 43650
rect 6414 43598 6466 43650
rect 7422 43598 7474 43650
rect 11118 43598 11170 43650
rect 17390 43598 17442 43650
rect 17614 43598 17666 43650
rect 17726 43598 17778 43650
rect 17838 43598 17890 43650
rect 18622 43598 18674 43650
rect 21646 43598 21698 43650
rect 26350 43598 26402 43650
rect 27134 43598 27186 43650
rect 29150 43598 29202 43650
rect 30942 43598 30994 43650
rect 31726 43598 31778 43650
rect 32062 43598 32114 43650
rect 33406 43598 33458 43650
rect 34638 43598 34690 43650
rect 37438 43598 37490 43650
rect 38782 43598 38834 43650
rect 39230 43598 39282 43650
rect 39454 43598 39506 43650
rect 39678 43598 39730 43650
rect 41582 43598 41634 43650
rect 2382 43486 2434 43538
rect 2494 43486 2546 43538
rect 2718 43486 2770 43538
rect 2942 43486 2994 43538
rect 4846 43486 4898 43538
rect 6974 43486 7026 43538
rect 8318 43486 8370 43538
rect 8766 43486 8818 43538
rect 9102 43486 9154 43538
rect 9998 43486 10050 43538
rect 10110 43486 10162 43538
rect 10894 43486 10946 43538
rect 12238 43486 12290 43538
rect 13022 43486 13074 43538
rect 13918 43486 13970 43538
rect 18510 43486 18562 43538
rect 20526 43486 20578 43538
rect 23438 43486 23490 43538
rect 23998 43486 24050 43538
rect 24670 43486 24722 43538
rect 25566 43486 25618 43538
rect 25678 43486 25730 43538
rect 25902 43486 25954 43538
rect 26574 43486 26626 43538
rect 28590 43486 28642 43538
rect 33182 43486 33234 43538
rect 33966 43486 34018 43538
rect 37326 43486 37378 43538
rect 41358 43486 41410 43538
rect 1822 43374 1874 43426
rect 2830 43374 2882 43426
rect 4062 43374 4114 43426
rect 4398 43374 4450 43426
rect 5854 43374 5906 43426
rect 6302 43374 6354 43426
rect 7870 43374 7922 43426
rect 10222 43374 10274 43426
rect 12350 43374 12402 43426
rect 12574 43374 12626 43426
rect 14478 43374 14530 43426
rect 23102 43374 23154 43426
rect 25342 43374 25394 43426
rect 32510 43374 32562 43426
rect 36766 43374 36818 43426
rect 41246 43374 41298 43426
rect 30718 43262 30770 43314
rect 31054 43262 31106 43314
rect 38670 43262 38722 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 24670 42926 24722 42978
rect 28366 42926 28418 42978
rect 13918 42814 13970 42866
rect 21758 42814 21810 42866
rect 25454 42814 25506 42866
rect 28254 42814 28306 42866
rect 30382 42814 30434 42866
rect 33854 42814 33906 42866
rect 34750 42814 34802 42866
rect 1822 42702 1874 42754
rect 7086 42702 7138 42754
rect 7646 42702 7698 42754
rect 8766 42702 8818 42754
rect 10782 42702 10834 42754
rect 13470 42702 13522 42754
rect 17614 42702 17666 42754
rect 18062 42702 18114 42754
rect 22542 42702 22594 42754
rect 25678 42702 25730 42754
rect 27022 42702 27074 42754
rect 29822 42702 29874 42754
rect 29934 42702 29986 42754
rect 30718 42702 30770 42754
rect 31166 42702 31218 42754
rect 33518 42702 33570 42754
rect 40126 42702 40178 42754
rect 40350 42702 40402 42754
rect 40686 42702 40738 42754
rect 41022 42702 41074 42754
rect 2046 42590 2098 42642
rect 2718 42590 2770 42642
rect 2830 42590 2882 42642
rect 9886 42590 9938 42642
rect 11342 42590 11394 42642
rect 24558 42590 24610 42642
rect 26238 42590 26290 42642
rect 30942 42590 30994 42642
rect 32958 42590 33010 42642
rect 3054 42478 3106 42530
rect 10894 42478 10946 42530
rect 21310 42478 21362 42530
rect 23102 42478 23154 42530
rect 23886 42478 23938 42530
rect 24334 42478 24386 42530
rect 24670 42478 24722 42530
rect 40686 42478 40738 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 3502 42142 3554 42194
rect 8878 42142 8930 42194
rect 16718 42142 16770 42194
rect 20974 42142 21026 42194
rect 29262 42142 29314 42194
rect 33182 42142 33234 42194
rect 35534 42142 35586 42194
rect 2270 42030 2322 42082
rect 6414 42030 6466 42082
rect 8430 42030 8482 42082
rect 11230 42030 11282 42082
rect 12126 42030 12178 42082
rect 16606 42030 16658 42082
rect 17838 42030 17890 42082
rect 17950 42030 18002 42082
rect 20750 42030 20802 42082
rect 26350 42030 26402 42082
rect 28590 42030 28642 42082
rect 30606 42030 30658 42082
rect 34526 42030 34578 42082
rect 35086 42030 35138 42082
rect 1822 41918 1874 41970
rect 2494 41918 2546 41970
rect 2718 41918 2770 41970
rect 2942 41918 2994 41970
rect 5294 41918 5346 41970
rect 7310 41918 7362 41970
rect 10558 41918 10610 41970
rect 12238 41918 12290 41970
rect 18398 41918 18450 41970
rect 18622 41918 18674 41970
rect 19966 41918 20018 41970
rect 20302 41918 20354 41970
rect 20526 41918 20578 41970
rect 20974 41918 21026 41970
rect 21982 41918 22034 41970
rect 22094 41918 22146 41970
rect 22206 41918 22258 41970
rect 22430 41918 22482 41970
rect 24782 41918 24834 41970
rect 25678 41918 25730 41970
rect 26238 41918 26290 41970
rect 26574 41918 26626 41970
rect 29710 41918 29762 41970
rect 30158 41918 30210 41970
rect 33966 41918 34018 41970
rect 35310 41918 35362 41970
rect 35870 41918 35922 41970
rect 40910 41918 40962 41970
rect 2606 41806 2658 41858
rect 4062 41806 4114 41858
rect 13358 41806 13410 41858
rect 18846 41806 18898 41858
rect 21534 41806 21586 41858
rect 22878 41806 22930 41858
rect 23214 41806 23266 41858
rect 25342 41806 25394 41858
rect 25902 41806 25954 41858
rect 26910 41806 26962 41858
rect 27582 41806 27634 41858
rect 32174 41806 32226 41858
rect 36318 41806 36370 41858
rect 40126 41806 40178 41858
rect 41694 41806 41746 41858
rect 43822 41806 43874 41858
rect 16718 41694 16770 41746
rect 17950 41694 18002 41746
rect 18958 41694 19010 41746
rect 34302 41694 34354 41746
rect 34638 41694 34690 41746
rect 35534 41694 35586 41746
rect 40014 41694 40066 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 12014 41358 12066 41410
rect 13918 41358 13970 41410
rect 14366 41358 14418 41410
rect 21758 41358 21810 41410
rect 21982 41358 22034 41410
rect 22094 41358 22146 41410
rect 27134 41358 27186 41410
rect 28030 41358 28082 41410
rect 30382 41358 30434 41410
rect 35422 41358 35474 41410
rect 7646 41246 7698 41298
rect 9550 41246 9602 41298
rect 18174 41246 18226 41298
rect 22878 41246 22930 41298
rect 25006 41246 25058 41298
rect 27806 41246 27858 41298
rect 28142 41246 28194 41298
rect 28590 41246 28642 41298
rect 30158 41246 30210 41298
rect 36094 41246 36146 41298
rect 37774 41246 37826 41298
rect 39902 41246 39954 41298
rect 1710 41134 1762 41186
rect 5854 41134 5906 41186
rect 9214 41134 9266 41186
rect 9326 41134 9378 41186
rect 11902 41134 11954 41186
rect 14142 41134 14194 41186
rect 17166 41134 17218 41186
rect 17614 41134 17666 41186
rect 19630 41134 19682 41186
rect 19966 41134 20018 41186
rect 20862 41134 20914 41186
rect 21422 41134 21474 41186
rect 21534 41134 21586 41186
rect 23214 41134 23266 41186
rect 24894 41134 24946 41186
rect 29150 41134 29202 41186
rect 29374 41134 29426 41186
rect 30494 41134 30546 41186
rect 31390 41134 31442 41186
rect 32958 41134 33010 41186
rect 33854 41134 33906 41186
rect 34862 41134 34914 41186
rect 35198 41134 35250 41186
rect 35422 41134 35474 41186
rect 36990 41134 37042 41186
rect 2046 41022 2098 41074
rect 2382 41022 2434 41074
rect 2718 41022 2770 41074
rect 6862 41022 6914 41074
rect 12126 41022 12178 41074
rect 13694 41022 13746 41074
rect 15710 41022 15762 41074
rect 19406 41022 19458 41074
rect 20526 41022 20578 41074
rect 23774 41022 23826 41074
rect 24782 41022 24834 41074
rect 31166 41022 31218 41074
rect 35982 41022 36034 41074
rect 7310 40910 7362 40962
rect 9662 40910 9714 40962
rect 14814 40910 14866 40962
rect 15150 40910 15202 40962
rect 19854 40910 19906 40962
rect 20638 40910 20690 40962
rect 27246 40910 27298 40962
rect 32958 40910 33010 40962
rect 35646 40910 35698 40962
rect 36206 40910 36258 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 12350 40574 12402 40626
rect 13134 40574 13186 40626
rect 16382 40574 16434 40626
rect 18174 40574 18226 40626
rect 19518 40574 19570 40626
rect 21086 40574 21138 40626
rect 22654 40574 22706 40626
rect 24110 40574 24162 40626
rect 25678 40574 25730 40626
rect 26686 40574 26738 40626
rect 27134 40574 27186 40626
rect 34078 40574 34130 40626
rect 34526 40574 34578 40626
rect 35758 40574 35810 40626
rect 36318 40574 36370 40626
rect 2046 40462 2098 40514
rect 4734 40462 4786 40514
rect 6190 40462 6242 40514
rect 9774 40462 9826 40514
rect 11790 40462 11842 40514
rect 15822 40462 15874 40514
rect 16158 40462 16210 40514
rect 17726 40462 17778 40514
rect 18622 40462 18674 40514
rect 34974 40462 35026 40514
rect 1710 40350 1762 40402
rect 2494 40350 2546 40402
rect 3390 40350 3442 40402
rect 5294 40350 5346 40402
rect 5742 40350 5794 40402
rect 8430 40350 8482 40402
rect 8654 40350 8706 40402
rect 9102 40350 9154 40402
rect 9998 40350 10050 40402
rect 12910 40350 12962 40402
rect 13582 40350 13634 40402
rect 14366 40350 14418 40402
rect 14814 40350 14866 40402
rect 15374 40350 15426 40402
rect 16606 40350 16658 40402
rect 17502 40350 17554 40402
rect 18846 40350 18898 40402
rect 19294 40350 19346 40402
rect 23102 40350 23154 40402
rect 26126 40350 26178 40402
rect 28254 40350 28306 40402
rect 28814 40350 28866 40402
rect 30494 40350 30546 40402
rect 30830 40350 30882 40402
rect 31166 40350 31218 40402
rect 35310 40350 35362 40402
rect 35422 40350 35474 40402
rect 35534 40350 35586 40402
rect 5406 40238 5458 40290
rect 8766 40238 8818 40290
rect 11342 40238 11394 40290
rect 12014 40238 12066 40290
rect 13022 40238 13074 40290
rect 18510 40238 18562 40290
rect 27806 40238 27858 40290
rect 29822 40238 29874 40290
rect 34638 40238 34690 40290
rect 36766 40238 36818 40290
rect 23774 40126 23826 40178
rect 24110 40126 24162 40178
rect 25342 40126 25394 40178
rect 25566 40126 25618 40178
rect 25678 40126 25730 40178
rect 26350 40126 26402 40178
rect 34302 40126 34354 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 7422 39790 7474 39842
rect 28702 39790 28754 39842
rect 30270 39790 30322 39842
rect 6078 39678 6130 39730
rect 11118 39678 11170 39730
rect 12686 39678 12738 39730
rect 22990 39678 23042 39730
rect 26686 39678 26738 39730
rect 29598 39678 29650 39730
rect 32286 39678 32338 39730
rect 3054 39566 3106 39618
rect 3950 39566 4002 39618
rect 5070 39566 5122 39618
rect 7982 39566 8034 39618
rect 8654 39566 8706 39618
rect 10670 39566 10722 39618
rect 10782 39566 10834 39618
rect 14142 39566 14194 39618
rect 14926 39566 14978 39618
rect 16382 39566 16434 39618
rect 17390 39566 17442 39618
rect 18734 39566 18786 39618
rect 21310 39566 21362 39618
rect 23326 39566 23378 39618
rect 27022 39566 27074 39618
rect 27806 39566 27858 39618
rect 28030 39566 28082 39618
rect 28254 39566 28306 39618
rect 30158 39566 30210 39618
rect 30718 39566 30770 39618
rect 30942 39566 30994 39618
rect 31390 39566 31442 39618
rect 31838 39566 31890 39618
rect 34078 39566 34130 39618
rect 34974 39566 35026 39618
rect 2830 39454 2882 39506
rect 3390 39454 3442 39506
rect 4958 39454 5010 39506
rect 7870 39454 7922 39506
rect 8766 39454 8818 39506
rect 18174 39454 18226 39506
rect 19630 39454 19682 39506
rect 22430 39454 22482 39506
rect 23886 39454 23938 39506
rect 25902 39454 25954 39506
rect 33854 39454 33906 39506
rect 34750 39454 34802 39506
rect 2942 39342 2994 39394
rect 3502 39342 3554 39394
rect 11566 39342 11618 39394
rect 14702 39342 14754 39394
rect 18062 39342 18114 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 3838 39006 3890 39058
rect 4286 39006 4338 39058
rect 5742 39006 5794 39058
rect 11790 39006 11842 39058
rect 13022 39006 13074 39058
rect 15262 39006 15314 39058
rect 19406 39006 19458 39058
rect 21982 39006 22034 39058
rect 22206 39006 22258 39058
rect 23774 39006 23826 39058
rect 24670 39006 24722 39058
rect 25118 39006 25170 39058
rect 27582 39006 27634 39058
rect 29598 39006 29650 39058
rect 2382 38894 2434 38946
rect 3502 38894 3554 38946
rect 5630 38894 5682 38946
rect 7086 38894 7138 38946
rect 15486 38894 15538 38946
rect 24222 38894 24274 38946
rect 26238 38894 26290 38946
rect 26798 38894 26850 38946
rect 28030 38894 28082 38946
rect 30942 38894 30994 38946
rect 32398 38894 32450 38946
rect 34302 38894 34354 38946
rect 35534 38894 35586 38946
rect 38222 38894 38274 38946
rect 2606 38782 2658 38834
rect 5182 38782 5234 38834
rect 6190 38782 6242 38834
rect 6526 38782 6578 38834
rect 7646 38782 7698 38834
rect 7870 38782 7922 38834
rect 12798 38782 12850 38834
rect 14030 38782 14082 38834
rect 14478 38782 14530 38834
rect 14814 38782 14866 38834
rect 15038 38782 15090 38834
rect 20974 38782 21026 38834
rect 21198 38782 21250 38834
rect 21310 38782 21362 38834
rect 21534 38782 21586 38834
rect 26014 38782 26066 38834
rect 26910 38782 26962 38834
rect 27134 38782 27186 38834
rect 28366 38782 28418 38834
rect 31278 38782 31330 38834
rect 31726 38782 31778 38834
rect 32510 38782 32562 38834
rect 34974 38782 35026 38834
rect 36878 38782 36930 38834
rect 37438 38782 37490 38834
rect 1822 38670 1874 38722
rect 7982 38670 8034 38722
rect 8542 38670 8594 38722
rect 12350 38670 12402 38722
rect 18062 38670 18114 38722
rect 18846 38670 18898 38722
rect 19966 38670 20018 38722
rect 20302 38670 20354 38722
rect 22766 38670 22818 38722
rect 23214 38670 23266 38722
rect 25566 38670 25618 38722
rect 26574 38670 26626 38722
rect 28142 38670 28194 38722
rect 28478 38670 28530 38722
rect 29038 38670 29090 38722
rect 33854 38670 33906 38722
rect 40350 38670 40402 38722
rect 7534 38558 7586 38610
rect 15374 38558 15426 38610
rect 25790 38558 25842 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 4958 38222 5010 38274
rect 13582 38222 13634 38274
rect 19070 38222 19122 38274
rect 20638 38222 20690 38274
rect 7422 38110 7474 38162
rect 11118 38110 11170 38162
rect 12238 38110 12290 38162
rect 15150 38110 15202 38162
rect 19630 38110 19682 38162
rect 27022 38110 27074 38162
rect 28366 38110 28418 38162
rect 29262 38110 29314 38162
rect 30046 38110 30098 38162
rect 32958 38110 33010 38162
rect 34302 38110 34354 38162
rect 37214 38110 37266 38162
rect 2494 37998 2546 38050
rect 3054 37998 3106 38050
rect 4062 37998 4114 38050
rect 4174 37998 4226 38050
rect 4734 37998 4786 38050
rect 5630 37998 5682 38050
rect 6526 37998 6578 38050
rect 7758 37998 7810 38050
rect 9550 37998 9602 38050
rect 9998 37998 10050 38050
rect 11454 37998 11506 38050
rect 11790 37998 11842 38050
rect 11902 37998 11954 38050
rect 12350 37998 12402 38050
rect 12798 37998 12850 38050
rect 14030 37998 14082 38050
rect 15038 37998 15090 38050
rect 15598 37998 15650 38050
rect 17278 37998 17330 38050
rect 17950 37998 18002 38050
rect 18398 37998 18450 38050
rect 18510 37998 18562 38050
rect 18734 37998 18786 38050
rect 18958 37998 19010 38050
rect 19966 37998 20018 38050
rect 20414 37998 20466 38050
rect 24110 37998 24162 38050
rect 26126 37998 26178 38050
rect 28254 37998 28306 38050
rect 28590 37998 28642 38050
rect 29822 37998 29874 38050
rect 30494 37998 30546 38050
rect 31838 37998 31890 38050
rect 33406 37998 33458 38050
rect 37774 37998 37826 38050
rect 37998 37998 38050 38050
rect 38222 37998 38274 38050
rect 1710 37886 1762 37938
rect 2606 37886 2658 37938
rect 4286 37886 4338 37938
rect 6974 37886 7026 37938
rect 10894 37886 10946 37938
rect 13470 37886 13522 37938
rect 14478 37886 14530 37938
rect 16942 37886 16994 37938
rect 17838 37886 17890 37938
rect 19742 37886 19794 37938
rect 22430 37886 22482 37938
rect 25230 37886 25282 37938
rect 26686 37886 26738 37938
rect 30606 37886 30658 37938
rect 32062 37886 32114 37938
rect 32174 37886 32226 37938
rect 38446 37886 38498 37938
rect 2046 37774 2098 37826
rect 2830 37774 2882 37826
rect 3614 37774 3666 37826
rect 6190 37774 6242 37826
rect 6862 37774 6914 37826
rect 9214 37774 9266 37826
rect 10670 37774 10722 37826
rect 11118 37774 11170 37826
rect 12126 37774 12178 37826
rect 13694 37774 13746 37826
rect 13918 37774 13970 37826
rect 15822 37774 15874 37826
rect 16382 37774 16434 37826
rect 17390 37774 17442 37826
rect 17614 37774 17666 37826
rect 21422 37774 21474 37826
rect 21870 37774 21922 37826
rect 22990 37774 23042 37826
rect 23438 37774 23490 37826
rect 23774 37774 23826 37826
rect 29710 37774 29762 37826
rect 33854 37774 33906 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2606 37438 2658 37490
rect 6302 37438 6354 37490
rect 8206 37438 8258 37490
rect 10558 37438 10610 37490
rect 12574 37438 12626 37490
rect 13022 37438 13074 37490
rect 15822 37438 15874 37490
rect 17950 37438 18002 37490
rect 24670 37438 24722 37490
rect 26686 37438 26738 37490
rect 28030 37438 28082 37490
rect 29038 37438 29090 37490
rect 29486 37438 29538 37490
rect 29710 37438 29762 37490
rect 32062 37438 32114 37490
rect 39566 37438 39618 37490
rect 39902 37438 39954 37490
rect 2046 37326 2098 37378
rect 2494 37326 2546 37378
rect 8766 37326 8818 37378
rect 9774 37326 9826 37378
rect 12126 37326 12178 37378
rect 16270 37326 16322 37378
rect 16494 37326 16546 37378
rect 18286 37326 18338 37378
rect 18398 37326 18450 37378
rect 19182 37326 19234 37378
rect 19406 37326 19458 37378
rect 23886 37326 23938 37378
rect 25790 37326 25842 37378
rect 26126 37326 26178 37378
rect 28254 37326 28306 37378
rect 29598 37326 29650 37378
rect 32286 37326 32338 37378
rect 35982 37326 36034 37378
rect 40350 37326 40402 37378
rect 1710 37214 1762 37266
rect 7758 37214 7810 37266
rect 8654 37214 8706 37266
rect 8990 37214 9042 37266
rect 9886 37214 9938 37266
rect 10110 37214 10162 37266
rect 11902 37214 11954 37266
rect 15374 37214 15426 37266
rect 15934 37214 15986 37266
rect 17614 37214 17666 37266
rect 18622 37214 18674 37266
rect 19070 37214 19122 37266
rect 20862 37214 20914 37266
rect 21086 37214 21138 37266
rect 21534 37214 21586 37266
rect 22766 37214 22818 37266
rect 24446 37214 24498 37266
rect 26462 37214 26514 37266
rect 27582 37214 27634 37266
rect 28366 37214 28418 37266
rect 29822 37214 29874 37266
rect 30046 37214 30098 37266
rect 31054 37214 31106 37266
rect 31278 37214 31330 37266
rect 31502 37214 31554 37266
rect 34302 37214 34354 37266
rect 34862 37214 34914 37266
rect 35310 37214 35362 37266
rect 3166 37102 3218 37154
rect 7422 37102 7474 37154
rect 9550 37102 9602 37154
rect 14926 37102 14978 37154
rect 25454 37102 25506 37154
rect 27806 37102 27858 37154
rect 31950 37102 32002 37154
rect 38110 37102 38162 37154
rect 2606 36990 2658 37042
rect 15150 36990 15202 37042
rect 16158 36990 16210 37042
rect 27134 36990 27186 37042
rect 27358 36990 27410 37042
rect 30494 36990 30546 37042
rect 40238 36990 40290 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 7198 36654 7250 36706
rect 14142 36654 14194 36706
rect 18174 36654 18226 36706
rect 18734 36654 18786 36706
rect 20078 36654 20130 36706
rect 3614 36542 3666 36594
rect 7086 36542 7138 36594
rect 8206 36542 8258 36594
rect 12910 36542 12962 36594
rect 17502 36542 17554 36594
rect 18846 36542 18898 36594
rect 27582 36542 27634 36594
rect 31726 36542 31778 36594
rect 33294 36542 33346 36594
rect 34638 36542 34690 36594
rect 36990 36542 37042 36594
rect 38894 36542 38946 36594
rect 2494 36430 2546 36482
rect 2718 36430 2770 36482
rect 3278 36430 3330 36482
rect 5742 36430 5794 36482
rect 8654 36430 8706 36482
rect 14366 36430 14418 36482
rect 18062 36430 18114 36482
rect 20414 36430 20466 36482
rect 20750 36430 20802 36482
rect 22542 36430 22594 36482
rect 24110 36430 24162 36482
rect 25790 36430 25842 36482
rect 26014 36430 26066 36482
rect 28702 36430 28754 36482
rect 29710 36430 29762 36482
rect 32174 36430 32226 36482
rect 32846 36430 32898 36482
rect 36318 36430 36370 36482
rect 39566 36430 39618 36482
rect 1934 36318 1986 36370
rect 3838 36318 3890 36370
rect 5966 36318 6018 36370
rect 6750 36318 6802 36370
rect 10446 36318 10498 36370
rect 13806 36318 13858 36370
rect 18286 36318 18338 36370
rect 20190 36318 20242 36370
rect 22878 36318 22930 36370
rect 23998 36318 24050 36370
rect 28366 36318 28418 36370
rect 35422 36318 35474 36370
rect 4286 36206 4338 36258
rect 4846 36206 4898 36258
rect 8990 36206 9042 36258
rect 14030 36206 14082 36258
rect 17838 36206 17890 36258
rect 19406 36206 19458 36258
rect 19742 36206 19794 36258
rect 20638 36206 20690 36258
rect 21534 36206 21586 36258
rect 21982 36206 22034 36258
rect 23886 36206 23938 36258
rect 28030 36206 28082 36258
rect 28478 36206 28530 36258
rect 29262 36206 29314 36258
rect 34078 36206 34130 36258
rect 37550 36206 37602 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 2494 35870 2546 35922
rect 2606 35870 2658 35922
rect 2830 35870 2882 35922
rect 3502 35870 3554 35922
rect 4622 35870 4674 35922
rect 5742 35870 5794 35922
rect 7646 35870 7698 35922
rect 9998 35870 10050 35922
rect 10222 35870 10274 35922
rect 10334 35870 10386 35922
rect 10670 35870 10722 35922
rect 11790 35870 11842 35922
rect 12014 35870 12066 35922
rect 12574 35870 12626 35922
rect 15038 35870 15090 35922
rect 18734 35870 18786 35922
rect 19742 35870 19794 35922
rect 20862 35870 20914 35922
rect 28702 35870 28754 35922
rect 29150 35870 29202 35922
rect 34750 35870 34802 35922
rect 37662 35870 37714 35922
rect 39342 35870 39394 35922
rect 2270 35758 2322 35810
rect 3726 35758 3778 35810
rect 14814 35758 14866 35810
rect 17726 35758 17778 35810
rect 19182 35758 19234 35810
rect 19966 35758 20018 35810
rect 20526 35758 20578 35810
rect 22878 35758 22930 35810
rect 23886 35758 23938 35810
rect 25454 35758 25506 35810
rect 27470 35758 27522 35810
rect 35646 35758 35698 35810
rect 37774 35758 37826 35810
rect 2718 35646 2770 35698
rect 3278 35646 3330 35698
rect 9662 35646 9714 35698
rect 12126 35646 12178 35698
rect 13918 35646 13970 35698
rect 14702 35646 14754 35698
rect 17614 35646 17666 35698
rect 18734 35646 18786 35698
rect 20078 35646 20130 35698
rect 20974 35646 21026 35698
rect 22990 35646 23042 35698
rect 23550 35646 23602 35698
rect 25230 35646 25282 35698
rect 27806 35646 27858 35698
rect 28254 35646 28306 35698
rect 33070 35646 33122 35698
rect 34750 35646 34802 35698
rect 38110 35646 38162 35698
rect 6302 35534 6354 35586
rect 8094 35534 8146 35586
rect 11566 35534 11618 35586
rect 13022 35534 13074 35586
rect 14366 35534 14418 35586
rect 15374 35534 15426 35586
rect 23214 35534 23266 35586
rect 25342 35534 25394 35586
rect 26686 35534 26738 35586
rect 27134 35534 27186 35586
rect 34190 35534 34242 35586
rect 36430 35534 36482 35586
rect 39790 35534 39842 35586
rect 3838 35422 3890 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 11566 35086 11618 35138
rect 12350 35086 12402 35138
rect 2830 34974 2882 35026
rect 9998 34974 10050 35026
rect 14814 34974 14866 35026
rect 17054 34974 17106 35026
rect 18734 34974 18786 35026
rect 26798 34974 26850 35026
rect 41918 34974 41970 35026
rect 2718 34862 2770 34914
rect 6190 34862 6242 34914
rect 6526 34862 6578 34914
rect 8094 34862 8146 34914
rect 8654 34862 8706 34914
rect 10446 34862 10498 34914
rect 10894 34862 10946 34914
rect 12238 34862 12290 34914
rect 12574 34862 12626 34914
rect 13470 34862 13522 34914
rect 14702 34862 14754 34914
rect 16494 34862 16546 34914
rect 16942 34862 16994 34914
rect 19294 34862 19346 34914
rect 19406 34862 19458 34914
rect 20190 34862 20242 34914
rect 20414 34862 20466 34914
rect 20750 34862 20802 34914
rect 22542 34862 22594 34914
rect 23774 34862 23826 34914
rect 25230 34862 25282 34914
rect 26574 34862 26626 34914
rect 27134 34862 27186 34914
rect 27582 34862 27634 34914
rect 27806 34862 27858 34914
rect 28254 34862 28306 34914
rect 29038 34862 29090 34914
rect 32398 34862 32450 34914
rect 32734 34862 32786 34914
rect 35086 34862 35138 34914
rect 36206 34862 36258 34914
rect 37326 34862 37378 34914
rect 39342 34862 39394 34914
rect 2270 34750 2322 34802
rect 2494 34750 2546 34802
rect 2830 34750 2882 34802
rect 5630 34750 5682 34802
rect 7646 34750 7698 34802
rect 11006 34750 11058 34802
rect 11118 34750 11170 34802
rect 13694 34750 13746 34802
rect 14926 34750 14978 34802
rect 15822 34750 15874 34802
rect 16830 34750 16882 34802
rect 18846 34750 18898 34802
rect 21646 34750 21698 34802
rect 23550 34750 23602 34802
rect 25342 34750 25394 34802
rect 25902 34750 25954 34802
rect 27022 34750 27074 34802
rect 29374 34750 29426 34802
rect 29822 34750 29874 34802
rect 33182 34750 33234 34802
rect 34526 34750 34578 34802
rect 36094 34750 36146 34802
rect 37438 34750 37490 34802
rect 39902 34750 39954 34802
rect 12014 34638 12066 34690
rect 12910 34638 12962 34690
rect 19070 34638 19122 34690
rect 20302 34638 20354 34690
rect 22766 34638 22818 34690
rect 26238 34638 26290 34690
rect 27694 34638 27746 34690
rect 28702 34638 28754 34690
rect 29262 34638 29314 34690
rect 30158 34638 30210 34690
rect 30942 34638 30994 34690
rect 31838 34638 31890 34690
rect 34638 34638 34690 34690
rect 37550 34638 37602 34690
rect 41470 34638 41522 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 1710 34302 1762 34354
rect 2494 34302 2546 34354
rect 3950 34302 4002 34354
rect 5406 34302 5458 34354
rect 7870 34302 7922 34354
rect 11566 34302 11618 34354
rect 13918 34302 13970 34354
rect 15822 34302 15874 34354
rect 17278 34302 17330 34354
rect 18062 34302 18114 34354
rect 18510 34302 18562 34354
rect 20078 34302 20130 34354
rect 39230 34302 39282 34354
rect 2046 34190 2098 34242
rect 10558 34190 10610 34242
rect 13134 34190 13186 34242
rect 14366 34190 14418 34242
rect 14814 34190 14866 34242
rect 15934 34190 15986 34242
rect 17502 34190 17554 34242
rect 19854 34190 19906 34242
rect 21870 34190 21922 34242
rect 23886 34190 23938 34242
rect 24222 34190 24274 34242
rect 25902 34190 25954 34242
rect 28030 34190 28082 34242
rect 28142 34190 28194 34242
rect 28254 34190 28306 34242
rect 33966 34190 34018 34242
rect 34862 34190 34914 34242
rect 37774 34190 37826 34242
rect 8542 34078 8594 34130
rect 9662 34078 9714 34130
rect 10670 34078 10722 34130
rect 12462 34078 12514 34130
rect 12910 34078 12962 34130
rect 14142 34078 14194 34130
rect 15262 34078 15314 34130
rect 16158 34078 16210 34130
rect 16718 34078 16770 34130
rect 17614 34078 17666 34130
rect 18398 34078 18450 34130
rect 18622 34078 18674 34130
rect 19070 34078 19122 34130
rect 20414 34078 20466 34130
rect 20974 34078 21026 34130
rect 21198 34078 21250 34130
rect 22206 34078 22258 34130
rect 22654 34078 22706 34130
rect 23550 34078 23602 34130
rect 23998 34078 24050 34130
rect 25342 34078 25394 34130
rect 25566 34078 25618 34130
rect 26238 34078 26290 34130
rect 30382 34078 30434 34130
rect 30830 34078 30882 34130
rect 31390 34078 31442 34130
rect 32510 34078 32562 34130
rect 34414 34078 34466 34130
rect 34750 34078 34802 34130
rect 36654 34078 36706 34130
rect 37102 34078 37154 34130
rect 38670 34078 38722 34130
rect 3502 33966 3554 34018
rect 5854 33966 5906 34018
rect 6638 33966 6690 34018
rect 7086 33966 7138 34018
rect 7422 33966 7474 34018
rect 8318 33966 8370 34018
rect 10110 33966 10162 34018
rect 11118 33966 11170 34018
rect 12014 33966 12066 34018
rect 19070 33966 19122 34018
rect 19518 33966 19570 34018
rect 8878 33854 8930 33906
rect 10558 33854 10610 33906
rect 11006 33854 11058 33906
rect 11678 33854 11730 33906
rect 24670 33966 24722 34018
rect 27246 33966 27298 34018
rect 28814 33966 28866 34018
rect 29262 33966 29314 34018
rect 29934 33966 29986 34018
rect 33630 33966 33682 34018
rect 39790 33966 39842 34018
rect 19630 33854 19682 33906
rect 27582 33854 27634 33906
rect 32398 33854 32450 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 13470 33518 13522 33570
rect 13918 33518 13970 33570
rect 14142 33518 14194 33570
rect 15038 33518 15090 33570
rect 18958 33518 19010 33570
rect 26798 33518 26850 33570
rect 8318 33406 8370 33458
rect 10110 33406 10162 33458
rect 14030 33406 14082 33458
rect 15038 33406 15090 33458
rect 15486 33406 15538 33458
rect 17166 33406 17218 33458
rect 20302 33406 20354 33458
rect 20750 33406 20802 33458
rect 23214 33406 23266 33458
rect 27918 33406 27970 33458
rect 33518 33406 33570 33458
rect 3278 33294 3330 33346
rect 4062 33294 4114 33346
rect 4286 33294 4338 33346
rect 4622 33294 4674 33346
rect 5070 33294 5122 33346
rect 5966 33294 6018 33346
rect 9214 33294 9266 33346
rect 9662 33294 9714 33346
rect 17614 33294 17666 33346
rect 18510 33294 18562 33346
rect 21534 33294 21586 33346
rect 23326 33294 23378 33346
rect 23774 33294 23826 33346
rect 25566 33294 25618 33346
rect 27806 33294 27858 33346
rect 28030 33294 28082 33346
rect 30382 33294 30434 33346
rect 32622 33294 32674 33346
rect 34750 33294 34802 33346
rect 35870 33294 35922 33346
rect 37102 33294 37154 33346
rect 39230 33294 39282 33346
rect 39566 33294 39618 33346
rect 1710 33182 1762 33234
rect 2494 33182 2546 33234
rect 2830 33182 2882 33234
rect 3726 33182 3778 33234
rect 4510 33182 4562 33234
rect 7422 33182 7474 33234
rect 8430 33182 8482 33234
rect 12126 33182 12178 33234
rect 12910 33182 12962 33234
rect 17166 33182 17218 33234
rect 19070 33182 19122 33234
rect 21982 33182 22034 33234
rect 25118 33182 25170 33234
rect 26350 33182 26402 33234
rect 28254 33182 28306 33234
rect 29262 33182 29314 33234
rect 34862 33182 34914 33234
rect 36318 33182 36370 33234
rect 38670 33182 38722 33234
rect 40126 33182 40178 33234
rect 2046 33070 2098 33122
rect 3838 33070 3890 33122
rect 12574 33070 12626 33122
rect 13694 33070 13746 33122
rect 14142 33070 14194 33122
rect 14590 33070 14642 33122
rect 16382 33070 16434 33122
rect 18286 33070 18338 33122
rect 18958 33070 19010 33122
rect 19518 33070 19570 33122
rect 22430 33070 22482 33122
rect 22878 33070 22930 33122
rect 23102 33070 23154 33122
rect 27694 33070 27746 33122
rect 30942 33070 30994 33122
rect 35310 33070 35362 33122
rect 37214 33070 37266 33122
rect 39006 33070 39058 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 5182 32734 5234 32786
rect 13470 32734 13522 32786
rect 19182 32734 19234 32786
rect 24670 32734 24722 32786
rect 28926 32734 28978 32786
rect 5406 32622 5458 32674
rect 14030 32622 14082 32674
rect 14366 32622 14418 32674
rect 16830 32622 16882 32674
rect 17950 32622 18002 32674
rect 21870 32622 21922 32674
rect 22318 32622 22370 32674
rect 28366 32622 28418 32674
rect 28478 32622 28530 32674
rect 33630 32622 33682 32674
rect 36206 32622 36258 32674
rect 2382 32510 2434 32562
rect 3278 32510 3330 32562
rect 3614 32510 3666 32562
rect 4958 32510 5010 32562
rect 6526 32510 6578 32562
rect 7310 32510 7362 32562
rect 8990 32510 9042 32562
rect 10334 32510 10386 32562
rect 12126 32510 12178 32562
rect 13246 32510 13298 32562
rect 17726 32510 17778 32562
rect 18846 32510 18898 32562
rect 21646 32510 21698 32562
rect 23662 32510 23714 32562
rect 25342 32510 25394 32562
rect 26350 32510 26402 32562
rect 27470 32510 27522 32562
rect 28142 32510 28194 32562
rect 33070 32510 33122 32562
rect 35086 32510 35138 32562
rect 38446 32510 38498 32562
rect 40014 32510 40066 32562
rect 8542 32398 8594 32450
rect 10670 32398 10722 32450
rect 12462 32398 12514 32450
rect 14814 32398 14866 32450
rect 15486 32398 15538 32450
rect 16494 32398 16546 32450
rect 18174 32398 18226 32450
rect 21422 32398 21474 32450
rect 23214 32398 23266 32450
rect 34862 32398 34914 32450
rect 37550 32398 37602 32450
rect 39566 32398 39618 32450
rect 26798 32286 26850 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 17390 31950 17442 32002
rect 2606 31838 2658 31890
rect 3502 31838 3554 31890
rect 18286 31838 18338 31890
rect 20414 31838 20466 31890
rect 24558 31838 24610 31890
rect 27134 31838 27186 31890
rect 29150 31838 29202 31890
rect 30494 31838 30546 31890
rect 3054 31726 3106 31778
rect 8990 31726 9042 31778
rect 9326 31726 9378 31778
rect 9662 31726 9714 31778
rect 11006 31726 11058 31778
rect 12798 31726 12850 31778
rect 13470 31726 13522 31778
rect 14030 31726 14082 31778
rect 15262 31726 15314 31778
rect 15822 31726 15874 31778
rect 16606 31726 16658 31778
rect 17054 31726 17106 31778
rect 17726 31726 17778 31778
rect 18510 31726 18562 31778
rect 19854 31726 19906 31778
rect 20190 31726 20242 31778
rect 20750 31726 20802 31778
rect 22430 31726 22482 31778
rect 22878 31726 22930 31778
rect 24894 31726 24946 31778
rect 26798 31726 26850 31778
rect 27358 31726 27410 31778
rect 33966 31726 34018 31778
rect 34302 31726 34354 31778
rect 36990 31726 37042 31778
rect 39118 31726 39170 31778
rect 11454 31614 11506 31666
rect 14590 31614 14642 31666
rect 14814 31614 14866 31666
rect 15038 31614 15090 31666
rect 16046 31614 16098 31666
rect 17950 31614 18002 31666
rect 24222 31614 24274 31666
rect 25230 31614 25282 31666
rect 27806 31614 27858 31666
rect 28030 31614 28082 31666
rect 33406 31614 33458 31666
rect 36094 31614 36146 31666
rect 37102 31614 37154 31666
rect 39678 31614 39730 31666
rect 3950 31502 4002 31554
rect 12910 31502 12962 31554
rect 14926 31502 14978 31554
rect 18958 31502 19010 31554
rect 19630 31502 19682 31554
rect 19742 31502 19794 31554
rect 20302 31502 20354 31554
rect 21422 31502 21474 31554
rect 29710 31502 29762 31554
rect 30942 31502 30994 31554
rect 32398 31502 32450 31554
rect 37214 31502 37266 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2270 31166 2322 31218
rect 9102 31166 9154 31218
rect 10894 31166 10946 31218
rect 13694 31166 13746 31218
rect 14142 31166 14194 31218
rect 14366 31166 14418 31218
rect 15150 31166 15202 31218
rect 15486 31166 15538 31218
rect 16270 31166 16322 31218
rect 17838 31166 17890 31218
rect 19070 31166 19122 31218
rect 20974 31166 21026 31218
rect 24222 31166 24274 31218
rect 24782 31166 24834 31218
rect 25790 31166 25842 31218
rect 26462 31166 26514 31218
rect 26686 31166 26738 31218
rect 27806 31166 27858 31218
rect 28478 31166 28530 31218
rect 28814 31166 28866 31218
rect 29038 31166 29090 31218
rect 33182 31166 33234 31218
rect 3054 31054 3106 31106
rect 4398 31054 4450 31106
rect 5630 31054 5682 31106
rect 12350 31054 12402 31106
rect 13918 31054 13970 31106
rect 17390 31054 17442 31106
rect 17614 31054 17666 31106
rect 18062 31054 18114 31106
rect 20078 31054 20130 31106
rect 20302 31054 20354 31106
rect 34302 31054 34354 31106
rect 35758 31054 35810 31106
rect 2158 30942 2210 30994
rect 3502 30942 3554 30994
rect 4286 30942 4338 30994
rect 6974 30942 7026 30994
rect 10110 30942 10162 30994
rect 11006 30942 11058 30994
rect 11902 30942 11954 30994
rect 14590 30942 14642 30994
rect 16158 30942 16210 30994
rect 18622 30942 18674 30994
rect 18734 30942 18786 30994
rect 18958 30942 19010 30994
rect 20638 30942 20690 30994
rect 26014 30942 26066 30994
rect 27246 30942 27298 30994
rect 27694 30942 27746 30994
rect 27918 30942 27970 30994
rect 29486 30942 29538 30994
rect 34862 30942 34914 30994
rect 36878 30942 36930 30994
rect 38222 30942 38274 30994
rect 3390 30830 3442 30882
rect 6302 30830 6354 30882
rect 7534 30830 7586 30882
rect 8654 30830 8706 30882
rect 14254 30830 14306 30882
rect 16830 30830 16882 30882
rect 18174 30830 18226 30882
rect 18846 30830 18898 30882
rect 19630 30830 19682 30882
rect 21422 30830 21474 30882
rect 21870 30830 21922 30882
rect 25342 30830 25394 30882
rect 26574 30830 26626 30882
rect 28926 30830 28978 30882
rect 37326 30830 37378 30882
rect 8654 30718 8706 30770
rect 9102 30718 9154 30770
rect 15150 30718 15202 30770
rect 15710 30718 15762 30770
rect 16270 30718 16322 30770
rect 20862 30718 20914 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 14366 30382 14418 30434
rect 14926 30382 14978 30434
rect 21870 30382 21922 30434
rect 26014 30382 26066 30434
rect 6526 30270 6578 30322
rect 9214 30270 9266 30322
rect 11790 30270 11842 30322
rect 14926 30270 14978 30322
rect 27022 30270 27074 30322
rect 30494 30270 30546 30322
rect 34414 30270 34466 30322
rect 36206 30270 36258 30322
rect 1710 30158 1762 30210
rect 4734 30158 4786 30210
rect 6190 30158 6242 30210
rect 6414 30158 6466 30210
rect 6862 30158 6914 30210
rect 7870 30158 7922 30210
rect 8430 30158 8482 30210
rect 9102 30158 9154 30210
rect 9886 30158 9938 30210
rect 12910 30158 12962 30210
rect 13582 30158 13634 30210
rect 14030 30158 14082 30210
rect 15486 30158 15538 30210
rect 17278 30158 17330 30210
rect 17502 30158 17554 30210
rect 18286 30158 18338 30210
rect 19294 30158 19346 30210
rect 19966 30158 20018 30210
rect 21534 30158 21586 30210
rect 21758 30158 21810 30210
rect 22430 30158 22482 30210
rect 23550 30158 23602 30210
rect 25006 30158 25058 30210
rect 25118 30158 25170 30210
rect 25454 30158 25506 30210
rect 26350 30158 26402 30210
rect 26574 30158 26626 30210
rect 28590 30158 28642 30210
rect 30942 30158 30994 30210
rect 31502 30158 31554 30210
rect 31950 30158 32002 30210
rect 34862 30158 34914 30210
rect 35870 30158 35922 30210
rect 2046 30046 2098 30098
rect 2382 30046 2434 30098
rect 4174 30046 4226 30098
rect 5070 30046 5122 30098
rect 7534 30046 7586 30098
rect 9662 30046 9714 30098
rect 11230 30046 11282 30098
rect 11678 30046 11730 30098
rect 12126 30046 12178 30098
rect 12574 30046 12626 30098
rect 12686 30046 12738 30098
rect 20414 30046 20466 30098
rect 21310 30046 21362 30098
rect 21982 30046 22034 30098
rect 22654 30046 22706 30098
rect 23102 30046 23154 30098
rect 23326 30046 23378 30098
rect 23998 30046 24050 30098
rect 24334 30046 24386 30098
rect 25230 30046 25282 30098
rect 25902 30046 25954 30098
rect 28142 30046 28194 30098
rect 2718 29934 2770 29986
rect 3166 29934 3218 29986
rect 4622 29934 4674 29986
rect 4958 29934 5010 29986
rect 5854 29934 5906 29986
rect 6638 29934 6690 29986
rect 10670 29934 10722 29986
rect 11566 29934 11618 29986
rect 11902 29934 11954 29986
rect 14478 29934 14530 29986
rect 26126 29934 26178 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 1822 29598 1874 29650
rect 6190 29598 6242 29650
rect 7086 29598 7138 29650
rect 11678 29598 11730 29650
rect 12686 29598 12738 29650
rect 15150 29598 15202 29650
rect 15710 29598 15762 29650
rect 2830 29486 2882 29538
rect 6414 29486 6466 29538
rect 7534 29486 7586 29538
rect 9774 29486 9826 29538
rect 2270 29374 2322 29426
rect 4622 29374 4674 29426
rect 5742 29374 5794 29426
rect 7982 29374 8034 29426
rect 8878 29374 8930 29426
rect 9662 29374 9714 29426
rect 10222 29374 10274 29426
rect 11006 29374 11058 29426
rect 12462 29374 12514 29426
rect 7646 29262 7698 29314
rect 12014 29262 12066 29314
rect 16158 29598 16210 29650
rect 18958 29598 19010 29650
rect 19518 29598 19570 29650
rect 20078 29598 20130 29650
rect 20862 29598 20914 29650
rect 23438 29598 23490 29650
rect 23774 29598 23826 29650
rect 23998 29598 24050 29650
rect 24222 29598 24274 29650
rect 25566 29598 25618 29650
rect 26014 29598 26066 29650
rect 27246 29598 27298 29650
rect 27806 29598 27858 29650
rect 35646 29598 35698 29650
rect 13694 29486 13746 29538
rect 14702 29486 14754 29538
rect 20414 29486 20466 29538
rect 27582 29486 27634 29538
rect 27918 29486 27970 29538
rect 28590 29486 28642 29538
rect 34190 29486 34242 29538
rect 37326 29486 37378 29538
rect 14366 29374 14418 29426
rect 14590 29374 14642 29426
rect 19742 29374 19794 29426
rect 19966 29374 20018 29426
rect 20190 29374 20242 29426
rect 21198 29374 21250 29426
rect 21758 29374 21810 29426
rect 22206 29374 22258 29426
rect 24334 29374 24386 29426
rect 28030 29374 28082 29426
rect 28366 29374 28418 29426
rect 28926 29374 28978 29426
rect 29598 29374 29650 29426
rect 35870 29374 35922 29426
rect 37886 29374 37938 29426
rect 22654 29262 22706 29314
rect 26686 29262 26738 29314
rect 10222 29150 10274 29202
rect 12686 29150 12738 29202
rect 13134 29150 13186 29202
rect 13358 29150 13410 29202
rect 13806 29150 13858 29202
rect 13918 29150 13970 29202
rect 15374 29150 15426 29202
rect 16158 29150 16210 29202
rect 25790 29150 25842 29202
rect 26126 29150 26178 29202
rect 29934 29150 29986 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21534 28814 21586 28866
rect 30158 28814 30210 28866
rect 2606 28702 2658 28754
rect 3838 28702 3890 28754
rect 6078 28702 6130 28754
rect 10670 28702 10722 28754
rect 11790 28702 11842 28754
rect 12126 28702 12178 28754
rect 12686 28702 12738 28754
rect 14478 28702 14530 28754
rect 15038 28702 15090 28754
rect 16606 28702 16658 28754
rect 20078 28702 20130 28754
rect 24558 28702 24610 28754
rect 26350 28702 26402 28754
rect 26910 28702 26962 28754
rect 27470 28702 27522 28754
rect 2270 28590 2322 28642
rect 2830 28590 2882 28642
rect 3950 28590 4002 28642
rect 6414 28590 6466 28642
rect 10110 28590 10162 28642
rect 10558 28590 10610 28642
rect 11230 28590 11282 28642
rect 15150 28590 15202 28642
rect 15262 28590 15314 28642
rect 16046 28590 16098 28642
rect 18510 28590 18562 28642
rect 18846 28590 18898 28642
rect 19294 28590 19346 28642
rect 20414 28590 20466 28642
rect 20750 28590 20802 28642
rect 21982 28590 22034 28642
rect 22542 28590 22594 28642
rect 23326 28590 23378 28642
rect 24670 28590 24722 28642
rect 25118 28590 25170 28642
rect 26014 28590 26066 28642
rect 28590 28590 28642 28642
rect 29150 28590 29202 28642
rect 29262 28590 29314 28642
rect 29486 28590 29538 28642
rect 29710 28590 29762 28642
rect 2494 28478 2546 28530
rect 3278 28478 3330 28530
rect 6974 28478 7026 28530
rect 10222 28478 10274 28530
rect 11006 28478 11058 28530
rect 14702 28478 14754 28530
rect 18734 28478 18786 28530
rect 21646 28478 21698 28530
rect 23438 28478 23490 28530
rect 24222 28478 24274 28530
rect 28254 28478 28306 28530
rect 28366 28478 28418 28530
rect 2718 28366 2770 28418
rect 3502 28366 3554 28418
rect 3726 28366 3778 28418
rect 6638 28366 6690 28418
rect 10782 28366 10834 28418
rect 14926 28366 14978 28418
rect 18286 28366 18338 28418
rect 20526 28366 20578 28418
rect 21534 28366 21586 28418
rect 28030 28366 28082 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 2046 28030 2098 28082
rect 4734 28030 4786 28082
rect 5182 28030 5234 28082
rect 7086 28030 7138 28082
rect 7982 28030 8034 28082
rect 8542 28030 8594 28082
rect 8654 28030 8706 28082
rect 8766 28030 8818 28082
rect 11454 28030 11506 28082
rect 13022 28030 13074 28082
rect 16270 28030 16322 28082
rect 16718 28030 16770 28082
rect 18174 28030 18226 28082
rect 22990 28030 23042 28082
rect 25454 28030 25506 28082
rect 25790 28030 25842 28082
rect 27022 28030 27074 28082
rect 29934 28030 29986 28082
rect 30830 28030 30882 28082
rect 4174 27918 4226 27970
rect 4958 27918 5010 27970
rect 5966 27918 6018 27970
rect 8990 27918 9042 27970
rect 12350 27918 12402 27970
rect 18398 27918 18450 27970
rect 19630 27918 19682 27970
rect 20638 27918 20690 27970
rect 20974 27918 21026 27970
rect 21646 27918 21698 27970
rect 27358 27918 27410 27970
rect 30270 27918 30322 27970
rect 1710 27806 1762 27858
rect 5518 27806 5570 27858
rect 5742 27806 5794 27858
rect 6638 27806 6690 27858
rect 6974 27806 7026 27858
rect 7758 27806 7810 27858
rect 8430 27806 8482 27858
rect 10558 27806 10610 27858
rect 12126 27806 12178 27858
rect 13694 27806 13746 27858
rect 14030 27806 14082 27858
rect 15486 27806 15538 27858
rect 15710 27806 15762 27858
rect 15822 27806 15874 27858
rect 16606 27806 16658 27858
rect 17726 27806 17778 27858
rect 17950 27806 18002 27858
rect 18734 27806 18786 27858
rect 19406 27806 19458 27858
rect 19966 27806 20018 27858
rect 21534 27806 21586 27858
rect 25678 27806 25730 27858
rect 25902 27806 25954 27858
rect 26462 27806 26514 27858
rect 27582 27806 27634 27858
rect 28142 27806 28194 27858
rect 29374 27806 29426 27858
rect 2494 27694 2546 27746
rect 5294 27694 5346 27746
rect 9998 27694 10050 27746
rect 24670 27694 24722 27746
rect 16718 27582 16770 27634
rect 17838 27582 17890 27634
rect 26686 27582 26738 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 17614 27246 17666 27298
rect 17838 27246 17890 27298
rect 24670 27246 24722 27298
rect 3726 27134 3778 27186
rect 4622 27134 4674 27186
rect 6414 27134 6466 27186
rect 8878 27134 8930 27186
rect 9214 27134 9266 27186
rect 10558 27134 10610 27186
rect 12574 27134 12626 27186
rect 14142 27134 14194 27186
rect 15262 27134 15314 27186
rect 17166 27134 17218 27186
rect 18062 27134 18114 27186
rect 18510 27134 18562 27186
rect 19406 27134 19458 27186
rect 20190 27134 20242 27186
rect 23774 27134 23826 27186
rect 27134 27134 27186 27186
rect 3950 27022 4002 27074
rect 4286 27022 4338 27074
rect 5854 27022 5906 27074
rect 9102 27022 9154 27074
rect 9774 27022 9826 27074
rect 14478 27022 14530 27074
rect 14702 27022 14754 27074
rect 15150 27022 15202 27074
rect 15710 27022 15762 27074
rect 16046 27022 16098 27074
rect 18622 27022 18674 27074
rect 24222 27022 24274 27074
rect 24446 27022 24498 27074
rect 25230 27022 25282 27074
rect 26014 27022 26066 27074
rect 3502 26910 3554 26962
rect 8094 26910 8146 26962
rect 10110 26910 10162 26962
rect 12126 26910 12178 26962
rect 13582 26910 13634 26962
rect 15374 26910 15426 26962
rect 15822 26910 15874 26962
rect 17614 26910 17666 26962
rect 18398 26910 18450 26962
rect 18846 26910 18898 26962
rect 25790 26910 25842 26962
rect 3726 26798 3778 26850
rect 9326 26798 9378 26850
rect 16606 26798 16658 26850
rect 21982 26798 22034 26850
rect 26574 26798 26626 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 9662 26462 9714 26514
rect 9774 26462 9826 26514
rect 10558 26462 10610 26514
rect 11006 26462 11058 26514
rect 12798 26462 12850 26514
rect 13246 26462 13298 26514
rect 13694 26462 13746 26514
rect 14142 26462 14194 26514
rect 14702 26462 14754 26514
rect 15598 26462 15650 26514
rect 17726 26462 17778 26514
rect 19518 26462 19570 26514
rect 20414 26462 20466 26514
rect 21758 26462 21810 26514
rect 26014 26462 26066 26514
rect 26574 26462 26626 26514
rect 7646 26350 7698 26402
rect 7870 26350 7922 26402
rect 15038 26350 15090 26402
rect 15710 26350 15762 26402
rect 17614 26350 17666 26402
rect 20862 26350 20914 26402
rect 5518 26238 5570 26290
rect 5966 26238 6018 26290
rect 7310 26238 7362 26290
rect 8206 26238 8258 26290
rect 9550 26238 9602 26290
rect 10110 26238 10162 26290
rect 11342 26238 11394 26290
rect 11902 26238 11954 26290
rect 12238 26238 12290 26290
rect 15486 26238 15538 26290
rect 15822 26238 15874 26290
rect 16046 26238 16098 26290
rect 17390 26238 17442 26290
rect 17838 26238 17890 26290
rect 17950 26238 18002 26290
rect 18510 26238 18562 26290
rect 21198 26238 21250 26290
rect 22206 26238 22258 26290
rect 8766 26126 8818 26178
rect 16830 26126 16882 26178
rect 19070 26126 19122 26178
rect 19966 26126 20018 26178
rect 22766 26126 22818 26178
rect 23214 26126 23266 26178
rect 25454 26126 25506 26178
rect 7086 26014 7138 26066
rect 7758 26014 7810 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 7310 25566 7362 25618
rect 8206 25566 8258 25618
rect 8542 25566 8594 25618
rect 14926 25566 14978 25618
rect 16494 25566 16546 25618
rect 17726 25566 17778 25618
rect 19966 25566 20018 25618
rect 27134 25566 27186 25618
rect 28254 25566 28306 25618
rect 29262 25566 29314 25618
rect 7646 25454 7698 25506
rect 8990 25454 9042 25506
rect 9438 25454 9490 25506
rect 9662 25454 9714 25506
rect 10222 25454 10274 25506
rect 10446 25454 10498 25506
rect 11006 25454 11058 25506
rect 11790 25454 11842 25506
rect 11902 25454 11954 25506
rect 12350 25454 12402 25506
rect 12910 25454 12962 25506
rect 14254 25454 14306 25506
rect 15262 25454 15314 25506
rect 16046 25454 16098 25506
rect 17390 25454 17442 25506
rect 18174 25454 18226 25506
rect 18846 25454 18898 25506
rect 19294 25454 19346 25506
rect 20078 25454 20130 25506
rect 21758 25454 21810 25506
rect 23662 25454 23714 25506
rect 25230 25454 25282 25506
rect 25566 25454 25618 25506
rect 27918 25454 27970 25506
rect 1710 25342 1762 25394
rect 2046 25342 2098 25394
rect 2494 25342 2546 25394
rect 6862 25342 6914 25394
rect 9550 25342 9602 25394
rect 10782 25342 10834 25394
rect 12574 25342 12626 25394
rect 14030 25342 14082 25394
rect 16382 25342 16434 25394
rect 17614 25342 17666 25394
rect 20414 25342 20466 25394
rect 22542 25342 22594 25394
rect 23550 25342 23602 25394
rect 9886 25230 9938 25282
rect 11342 25230 11394 25282
rect 12014 25230 12066 25282
rect 12798 25230 12850 25282
rect 13694 25230 13746 25282
rect 15262 25230 15314 25282
rect 18622 25230 18674 25282
rect 21534 25230 21586 25282
rect 21870 25230 21922 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 11230 24894 11282 24946
rect 11678 24894 11730 24946
rect 16718 24894 16770 24946
rect 17614 24894 17666 24946
rect 22990 24894 23042 24946
rect 16046 24782 16098 24834
rect 19294 24782 19346 24834
rect 20414 24782 20466 24834
rect 22430 24782 22482 24834
rect 24222 24782 24274 24834
rect 13022 24670 13074 24722
rect 13358 24670 13410 24722
rect 13582 24670 13634 24722
rect 13918 24670 13970 24722
rect 16494 24670 16546 24722
rect 17838 24670 17890 24722
rect 21086 24670 21138 24722
rect 21982 24670 22034 24722
rect 24446 24670 24498 24722
rect 25790 24670 25842 24722
rect 19182 24558 19234 24610
rect 25342 24558 25394 24610
rect 26238 24558 26290 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 20750 24110 20802 24162
rect 11678 23998 11730 24050
rect 12462 23998 12514 24050
rect 14030 23998 14082 24050
rect 15150 23998 15202 24050
rect 16158 23998 16210 24050
rect 19742 23998 19794 24050
rect 21534 23998 21586 24050
rect 23438 23998 23490 24050
rect 24222 23998 24274 24050
rect 25230 23998 25282 24050
rect 25790 23998 25842 24050
rect 12910 23886 12962 23938
rect 14702 23886 14754 23938
rect 15598 23886 15650 23938
rect 16382 23886 16434 23938
rect 17950 23886 18002 23938
rect 19966 23886 20018 23938
rect 20190 23886 20242 23938
rect 20302 23886 20354 23938
rect 21982 23886 22034 23938
rect 22318 23886 22370 23938
rect 23774 23886 23826 23938
rect 24782 23886 24834 23938
rect 1710 23774 1762 23826
rect 2046 23774 2098 23826
rect 16942 23774 16994 23826
rect 18174 23774 18226 23826
rect 21310 23774 21362 23826
rect 2494 23662 2546 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 15150 23326 15202 23378
rect 15598 23326 15650 23378
rect 15934 23326 15986 23378
rect 16158 23326 16210 23378
rect 16606 23326 16658 23378
rect 19070 23326 19122 23378
rect 21086 23326 21138 23378
rect 21646 23326 21698 23378
rect 22990 23326 23042 23378
rect 25454 23326 25506 23378
rect 15822 23214 15874 23266
rect 19182 23214 19234 23266
rect 21310 23214 21362 23266
rect 22206 23214 22258 23266
rect 17614 22990 17666 23042
rect 19070 22878 19122 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 1710 22206 1762 22258
rect 2046 22206 2098 22258
rect 2494 22094 2546 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 2046 20638 2098 20690
rect 1710 20526 1762 20578
rect 2494 20526 2546 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 2046 18622 2098 18674
rect 1710 18398 1762 18450
rect 2494 18286 2546 18338
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 2046 17054 2098 17106
rect 1710 16830 1762 16882
rect 2494 16830 2546 16882
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 2046 15486 2098 15538
rect 1710 15262 1762 15314
rect 2494 15150 2546 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 1710 12798 1762 12850
rect 2046 12798 2098 12850
rect 2494 12798 2546 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 1710 11230 1762 11282
rect 2046 11230 2098 11282
rect 2494 11118 2546 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 1710 9662 1762 9714
rect 2046 9662 2098 9714
rect 2494 9550 2546 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 1710 8094 1762 8146
rect 2046 8094 2098 8146
rect 2494 7982 2546 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 1710 5854 1762 5906
rect 2158 5742 2210 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 1822 5182 1874 5234
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 2046 4510 2098 4562
rect 1710 4286 1762 4338
rect 2494 4174 2546 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 2270 3614 2322 3666
rect 1710 3390 1762 3442
rect 2718 3390 2770 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 2912 59200 3024 60000
rect 5152 59200 5264 60000
rect 7392 59200 7504 60000
rect 9632 59200 9744 60000
rect 11872 59200 11984 60000
rect 14112 59200 14224 60000
rect 16352 59200 16464 60000
rect 18592 59200 18704 60000
rect 20832 59200 20944 60000
rect 23072 59200 23184 60000
rect 25312 59200 25424 60000
rect 27552 59200 27664 60000
rect 29792 59200 29904 60000
rect 32032 59200 32144 60000
rect 34272 59200 34384 60000
rect 36512 59200 36624 60000
rect 38752 59200 38864 60000
rect 40992 59200 41104 60000
rect 43232 59200 43344 60000
rect 45472 59200 45584 60000
rect 47712 59200 47824 60000
rect 49952 59200 50064 60000
rect 52192 59200 52304 60000
rect 54432 59200 54544 60000
rect 56672 59200 56784 60000
rect 2156 57652 2212 57662
rect 2044 56194 2100 56206
rect 2044 56142 2046 56194
rect 2098 56142 2100 56194
rect 1708 56082 1764 56094
rect 1708 56030 1710 56082
rect 1762 56030 1764 56082
rect 1708 55860 1764 56030
rect 1708 55794 1764 55804
rect 2044 55468 2100 56142
rect 1932 55412 2100 55468
rect 2156 56084 2212 57596
rect 1596 54628 1652 54638
rect 1484 44884 1540 44894
rect 924 42308 980 42318
rect 924 28756 980 42252
rect 1036 39620 1092 39630
rect 1036 32900 1092 39564
rect 1372 36260 1428 36270
rect 1036 32834 1092 32844
rect 1148 35700 1204 35710
rect 924 28690 980 28700
rect 1036 32452 1092 32462
rect 1036 5908 1092 32396
rect 1148 23492 1204 35644
rect 1148 23426 1204 23436
rect 1372 15764 1428 36204
rect 1484 28308 1540 44828
rect 1596 36484 1652 54572
rect 1708 54514 1764 54526
rect 1708 54462 1710 54514
rect 1762 54462 1764 54514
rect 1708 54068 1764 54462
rect 1708 54002 1764 54012
rect 1708 52946 1764 52958
rect 1708 52894 1710 52946
rect 1762 52894 1764 52946
rect 1708 52836 1764 52894
rect 1708 52276 1764 52780
rect 1708 52210 1764 52220
rect 1820 51378 1876 51390
rect 1820 51326 1822 51378
rect 1874 51326 1876 51378
rect 1820 51268 1876 51326
rect 1708 50708 1764 50718
rect 1708 50614 1764 50652
rect 1708 50484 1764 50494
rect 1820 50484 1876 51212
rect 1764 50428 1876 50484
rect 1708 50418 1764 50428
rect 1932 49812 1988 55412
rect 2156 55410 2212 56028
rect 2156 55358 2158 55410
rect 2210 55358 2212 55410
rect 2156 55346 2212 55358
rect 2380 56194 2436 56206
rect 2380 56142 2382 56194
rect 2434 56142 2436 56194
rect 2044 54628 2100 54638
rect 2044 54534 2100 54572
rect 2044 53060 2100 53070
rect 2044 53058 2324 53060
rect 2044 53006 2046 53058
rect 2098 53006 2324 53058
rect 2044 53004 2324 53006
rect 2044 52994 2100 53004
rect 2268 52722 2324 53004
rect 2268 52670 2270 52722
rect 2322 52670 2324 52722
rect 2268 52658 2324 52670
rect 2044 51492 2100 51502
rect 2044 51398 2100 51436
rect 2044 50708 2100 50718
rect 2100 50652 2324 50708
rect 2044 50642 2100 50652
rect 2268 50036 2324 50652
rect 2268 49970 2324 49980
rect 1932 49756 2324 49812
rect 1708 49700 1764 49710
rect 1708 49698 2212 49700
rect 1708 49646 1710 49698
rect 1762 49646 2212 49698
rect 1708 49644 2212 49646
rect 1708 49634 1764 49644
rect 1708 48914 1764 48926
rect 1708 48862 1710 48914
rect 1762 48862 1764 48914
rect 1708 48692 1764 48862
rect 2044 48804 2100 48814
rect 1708 48626 1764 48636
rect 1820 48802 2100 48804
rect 1820 48750 2046 48802
rect 2098 48750 2100 48802
rect 1820 48748 2100 48750
rect 1708 46900 1764 46910
rect 1708 46786 1764 46844
rect 1708 46734 1710 46786
rect 1762 46734 1764 46786
rect 1708 46722 1764 46734
rect 1708 45778 1764 45790
rect 1708 45726 1710 45778
rect 1762 45726 1764 45778
rect 1708 45332 1764 45726
rect 1708 45108 1764 45276
rect 1708 45042 1764 45052
rect 1820 43652 1876 48748
rect 2044 48738 2100 48748
rect 2156 47684 2212 49644
rect 2156 47458 2212 47628
rect 2156 47406 2158 47458
rect 2210 47406 2212 47458
rect 2156 47394 2212 47406
rect 2044 46788 2100 46798
rect 1820 43586 1876 43596
rect 1932 46786 2100 46788
rect 1932 46734 2046 46786
rect 2098 46734 2100 46786
rect 1932 46732 2100 46734
rect 1820 43426 1876 43438
rect 1820 43374 1822 43426
rect 1874 43374 1876 43426
rect 1820 43316 1876 43374
rect 1820 42754 1876 43260
rect 1820 42702 1822 42754
rect 1874 42702 1876 42754
rect 1820 42690 1876 42702
rect 1820 41972 1876 41982
rect 1708 41970 1876 41972
rect 1708 41918 1822 41970
rect 1874 41918 1876 41970
rect 1708 41916 1876 41918
rect 1708 41524 1764 41916
rect 1820 41906 1876 41916
rect 1708 41186 1764 41468
rect 1708 41134 1710 41186
rect 1762 41134 1764 41186
rect 1708 41122 1764 41134
rect 1708 40402 1764 40414
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 40292 1764 40350
rect 1708 39732 1764 40236
rect 1708 39666 1764 39676
rect 1932 39396 1988 46732
rect 2044 46722 2100 46732
rect 2044 45668 2100 45678
rect 2044 45666 2212 45668
rect 2044 45614 2046 45666
rect 2098 45614 2212 45666
rect 2044 45612 2212 45614
rect 2044 45602 2100 45612
rect 2044 43540 2100 43550
rect 2044 42642 2100 43484
rect 2044 42590 2046 42642
rect 2098 42590 2100 42642
rect 2044 42578 2100 42590
rect 2156 42532 2212 45612
rect 2268 44548 2324 49756
rect 2268 44482 2324 44492
rect 2380 43538 2436 56142
rect 2604 56084 2660 56094
rect 2604 55990 2660 56028
rect 2492 54402 2548 54414
rect 2492 54350 2494 54402
rect 2546 54350 2548 54402
rect 2492 54068 2548 54350
rect 2492 54002 2548 54012
rect 2940 53844 2996 59200
rect 5068 56308 5124 56318
rect 5180 56308 5236 59200
rect 7420 56308 7476 59200
rect 7644 56308 7700 56318
rect 5068 56306 5572 56308
rect 5068 56254 5070 56306
rect 5122 56254 5572 56306
rect 5068 56252 5572 56254
rect 5068 56242 5124 56252
rect 5516 56194 5572 56252
rect 7420 56306 7700 56308
rect 7420 56254 7422 56306
rect 7474 56254 7646 56306
rect 7698 56254 7700 56306
rect 7420 56252 7700 56254
rect 7420 56242 7476 56252
rect 7644 56242 7700 56252
rect 9660 56308 9716 59200
rect 9884 56308 9940 56318
rect 9660 56306 9940 56308
rect 9660 56254 9662 56306
rect 9714 56254 9886 56306
rect 9938 56254 9940 56306
rect 9660 56252 9940 56254
rect 9660 56242 9716 56252
rect 9884 56242 9940 56252
rect 11900 56308 11956 59200
rect 14140 56420 14196 59200
rect 14140 56364 14644 56420
rect 12124 56308 12180 56318
rect 11900 56306 12180 56308
rect 11900 56254 11902 56306
rect 11954 56254 12126 56306
rect 12178 56254 12180 56306
rect 11900 56252 12180 56254
rect 11900 56242 11956 56252
rect 12124 56242 12180 56252
rect 14140 56306 14196 56364
rect 14140 56254 14142 56306
rect 14194 56254 14196 56306
rect 14140 56242 14196 56254
rect 5516 56142 5518 56194
rect 5570 56142 5572 56194
rect 5516 56130 5572 56142
rect 5852 56194 5908 56206
rect 5852 56142 5854 56194
rect 5906 56142 5908 56194
rect 3164 55970 3220 55982
rect 3164 55918 3166 55970
rect 3218 55918 3220 55970
rect 3164 55860 3220 55918
rect 3164 55794 3220 55804
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 5852 55188 5908 56142
rect 7980 56194 8036 56206
rect 7980 56142 7982 56194
rect 8034 56142 8036 56194
rect 7980 55468 8036 56142
rect 10220 56194 10276 56206
rect 10220 56142 10222 56194
rect 10274 56142 10276 56194
rect 10220 55468 10276 56142
rect 12460 56194 12516 56206
rect 12460 56142 12462 56194
rect 12514 56142 12516 56194
rect 12460 55468 12516 56142
rect 14364 56194 14420 56206
rect 14364 56142 14366 56194
rect 14418 56142 14420 56194
rect 14364 55468 14420 56142
rect 14588 56082 14644 56364
rect 16380 56308 16436 59200
rect 16492 56308 16548 56318
rect 16940 56308 16996 56318
rect 16380 56306 16996 56308
rect 16380 56254 16494 56306
rect 16546 56254 16942 56306
rect 16994 56254 16996 56306
rect 16380 56252 16996 56254
rect 16492 56242 16548 56252
rect 16940 56242 16996 56252
rect 18620 56308 18676 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 18844 56308 18900 56318
rect 18620 56306 18900 56308
rect 18620 56254 18622 56306
rect 18674 56254 18846 56306
rect 18898 56254 18900 56306
rect 18620 56252 18900 56254
rect 18620 56242 18676 56252
rect 18844 56242 18900 56252
rect 20300 56308 20356 56318
rect 20860 56308 20916 59200
rect 20300 56306 20916 56308
rect 20300 56254 20302 56306
rect 20354 56254 20916 56306
rect 20300 56252 20916 56254
rect 20300 56242 20356 56252
rect 17276 56196 17332 56206
rect 17276 56194 17556 56196
rect 17276 56142 17278 56194
rect 17330 56142 17556 56194
rect 17276 56140 17556 56142
rect 17276 56130 17332 56140
rect 14588 56030 14590 56082
rect 14642 56030 14644 56082
rect 14588 56018 14644 56030
rect 7980 55412 8260 55468
rect 10220 55412 10500 55468
rect 5852 55122 5908 55132
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 2940 53778 2996 53788
rect 5628 53844 5684 53854
rect 2492 52836 2548 52846
rect 2492 52742 2548 52780
rect 2604 52722 2660 52734
rect 2604 52670 2606 52722
rect 2658 52670 2660 52722
rect 2492 51268 2548 51278
rect 2492 51174 2548 51212
rect 2492 48802 2548 48814
rect 2492 48750 2494 48802
rect 2546 48750 2548 48802
rect 2492 48692 2548 48750
rect 2492 48626 2548 48636
rect 2492 46900 2548 46910
rect 2492 46806 2548 46844
rect 2492 45666 2548 45678
rect 2492 45614 2494 45666
rect 2546 45614 2548 45666
rect 2492 45332 2548 45614
rect 2492 45266 2548 45276
rect 2604 45330 2660 52670
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 3836 51940 3892 51950
rect 2716 51492 2772 51502
rect 2772 51436 2884 51492
rect 2716 51426 2772 51436
rect 2716 50036 2772 50046
rect 2716 48468 2772 49980
rect 2716 48402 2772 48412
rect 2716 47460 2772 47470
rect 2716 47366 2772 47404
rect 2828 46116 2884 51436
rect 3836 50706 3892 51884
rect 5628 51492 5684 53788
rect 7980 53060 8036 53070
rect 7980 52966 8036 53004
rect 5628 51426 5684 51436
rect 5852 52834 5908 52846
rect 5852 52782 5854 52834
rect 5906 52782 5908 52834
rect 4396 51380 4452 51390
rect 4396 51286 4452 51324
rect 5180 51380 5236 51390
rect 5068 51268 5124 51278
rect 5068 51174 5124 51212
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 5068 50708 5124 50718
rect 5180 50708 5236 51324
rect 5852 50820 5908 52782
rect 7644 51380 7700 51390
rect 7644 51286 7700 51324
rect 7196 51268 7252 51278
rect 5852 50754 5908 50764
rect 7084 51266 7252 51268
rect 7084 51214 7198 51266
rect 7250 51214 7252 51266
rect 7084 51212 7252 51214
rect 7084 50708 7140 51212
rect 7196 51202 7252 51212
rect 7308 50820 7364 50830
rect 3836 50654 3838 50706
rect 3890 50654 3892 50706
rect 3836 50642 3892 50654
rect 4620 50706 5236 50708
rect 4620 50654 5070 50706
rect 5122 50654 5236 50706
rect 4620 50652 5236 50654
rect 6748 50706 7140 50708
rect 6748 50654 7086 50706
rect 7138 50654 7140 50706
rect 6748 50652 7140 50654
rect 4620 50594 4676 50652
rect 4620 50542 4622 50594
rect 4674 50542 4676 50594
rect 3836 49924 3892 49934
rect 3836 49830 3892 49868
rect 4620 49810 4676 50542
rect 5068 50034 5124 50652
rect 6748 50428 6804 50652
rect 5068 49982 5070 50034
rect 5122 49982 5124 50034
rect 5068 49970 5124 49982
rect 6524 50372 6804 50428
rect 4620 49758 4622 49810
rect 4674 49758 4676 49810
rect 4620 49746 4676 49758
rect 6524 49810 6580 50372
rect 6524 49758 6526 49810
rect 6578 49758 6580 49810
rect 6524 49746 6580 49758
rect 6412 49698 6468 49710
rect 6412 49646 6414 49698
rect 6466 49646 6468 49698
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 3052 48468 3108 48478
rect 3052 47570 3108 48412
rect 3500 48468 3556 48478
rect 3500 48374 3556 48412
rect 4060 48130 4116 48142
rect 4060 48078 4062 48130
rect 4114 48078 4116 48130
rect 3276 47684 3332 47694
rect 3276 47590 3332 47628
rect 3052 47518 3054 47570
rect 3106 47518 3108 47570
rect 2940 46788 2996 46798
rect 3052 46788 3108 47518
rect 3948 47460 4004 47470
rect 2940 46786 3108 46788
rect 2940 46734 2942 46786
rect 2994 46734 3108 46786
rect 2940 46732 3108 46734
rect 3612 47234 3668 47246
rect 3612 47182 3614 47234
rect 3666 47182 3668 47234
rect 2940 46722 2996 46732
rect 3052 46452 3108 46462
rect 3052 46450 3332 46452
rect 3052 46398 3054 46450
rect 3106 46398 3332 46450
rect 3052 46396 3332 46398
rect 3052 46386 3108 46396
rect 2828 46060 3220 46116
rect 2604 45278 2606 45330
rect 2658 45278 2660 45330
rect 2604 45266 2660 45278
rect 3164 45330 3220 46060
rect 3164 45278 3166 45330
rect 3218 45278 3220 45330
rect 3164 45266 3220 45278
rect 2380 43486 2382 43538
rect 2434 43486 2436 43538
rect 2380 43474 2436 43486
rect 2492 45108 2548 45118
rect 3052 45108 3108 45118
rect 2492 45106 3108 45108
rect 2492 45054 2494 45106
rect 2546 45054 3054 45106
rect 3106 45054 3108 45106
rect 2492 45052 3108 45054
rect 3276 45108 3332 46396
rect 3276 45052 3556 45108
rect 2492 43538 2548 45052
rect 3052 45042 3108 45052
rect 2604 44884 2660 44894
rect 3164 44884 3220 44894
rect 2604 44882 3108 44884
rect 2604 44830 2606 44882
rect 2658 44830 3108 44882
rect 2604 44828 3108 44830
rect 2604 44818 2660 44828
rect 2492 43486 2494 43538
rect 2546 43486 2548 43538
rect 2156 42476 2436 42532
rect 2268 42084 2324 42094
rect 2268 41990 2324 42028
rect 2044 41972 2100 41982
rect 2044 41074 2100 41916
rect 2380 41300 2436 42476
rect 2044 41022 2046 41074
rect 2098 41022 2100 41074
rect 2044 41010 2100 41022
rect 2268 41244 2436 41300
rect 2492 41970 2548 43486
rect 2716 43540 2772 43550
rect 2716 43446 2772 43484
rect 2940 43538 2996 43550
rect 2940 43486 2942 43538
rect 2994 43486 2996 43538
rect 2828 43426 2884 43438
rect 2828 43374 2830 43426
rect 2882 43374 2884 43426
rect 2716 42644 2772 42654
rect 2716 42550 2772 42588
rect 2828 42642 2884 43374
rect 2828 42590 2830 42642
rect 2882 42590 2884 42642
rect 2828 42578 2884 42590
rect 2492 41918 2494 41970
rect 2546 41918 2548 41970
rect 2044 40514 2100 40526
rect 2044 40462 2046 40514
rect 2098 40462 2100 40514
rect 2044 39620 2100 40462
rect 2044 39554 2100 39564
rect 1932 39340 2212 39396
rect 1820 38722 1876 38734
rect 1820 38670 1822 38722
rect 1874 38670 1876 38722
rect 1820 38668 1876 38670
rect 1708 38612 1876 38668
rect 1708 37940 1764 38612
rect 1708 37846 1764 37884
rect 2044 37828 2100 37838
rect 2044 37734 2100 37772
rect 2044 37380 2100 37390
rect 1820 37378 2100 37380
rect 1820 37326 2046 37378
rect 2098 37326 2100 37378
rect 1820 37324 2100 37326
rect 1596 36418 1652 36428
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 37156 1764 37214
rect 1708 36148 1764 37100
rect 1708 36082 1764 36092
rect 1484 28242 1540 28252
rect 1596 34468 1652 34478
rect 1372 15698 1428 15708
rect 1036 5842 1092 5852
rect 1596 4564 1652 34412
rect 1708 34356 1764 34366
rect 1708 34262 1764 34300
rect 1708 33236 1764 33246
rect 1708 32564 1764 33180
rect 1708 32498 1764 32508
rect 1820 31108 1876 37324
rect 2044 37314 2100 37324
rect 2044 36596 2100 36606
rect 1932 36372 1988 36382
rect 1932 36278 1988 36316
rect 1820 31042 1876 31052
rect 1932 36036 1988 36046
rect 1708 30772 1764 30782
rect 1708 30212 1764 30716
rect 1708 30210 1876 30212
rect 1708 30158 1710 30210
rect 1762 30158 1876 30210
rect 1708 30156 1876 30158
rect 1708 30146 1764 30156
rect 1820 29650 1876 30156
rect 1820 29598 1822 29650
rect 1874 29598 1876 29650
rect 1820 29586 1876 29598
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27748 1764 27806
rect 1708 27188 1764 27692
rect 1708 27122 1764 27132
rect 1708 25396 1764 25406
rect 1932 25396 1988 35980
rect 2044 35252 2100 36540
rect 2156 35812 2212 39340
rect 2268 39172 2324 41244
rect 2492 41188 2548 41918
rect 2716 41972 2772 41982
rect 2716 41878 2772 41916
rect 2940 41972 2996 43486
rect 3052 42756 3108 44828
rect 3164 44790 3220 44828
rect 3500 43650 3556 45052
rect 3500 43598 3502 43650
rect 3554 43598 3556 43650
rect 3052 42700 3332 42756
rect 3052 42532 3108 42542
rect 3052 42438 3108 42476
rect 2940 41970 3220 41972
rect 2940 41918 2942 41970
rect 2994 41918 3220 41970
rect 2940 41916 3220 41918
rect 2940 41906 2996 41916
rect 2604 41858 2660 41870
rect 2604 41806 2606 41858
rect 2658 41806 2660 41858
rect 2604 41300 2660 41806
rect 2604 41244 2996 41300
rect 2492 41132 2772 41188
rect 2380 41074 2436 41086
rect 2380 41022 2382 41074
rect 2434 41022 2436 41074
rect 2380 39620 2436 41022
rect 2716 41074 2772 41132
rect 2716 41022 2718 41074
rect 2770 41022 2772 41074
rect 2716 41010 2772 41022
rect 2492 40402 2548 40414
rect 2492 40350 2494 40402
rect 2546 40350 2548 40402
rect 2492 40292 2548 40350
rect 2492 40226 2548 40236
rect 2828 40292 2884 40302
rect 2380 39564 2660 39620
rect 2268 39116 2548 39172
rect 2380 38946 2436 38958
rect 2380 38894 2382 38946
rect 2434 38894 2436 38946
rect 2380 38052 2436 38894
rect 2492 38668 2548 39116
rect 2604 39060 2660 39564
rect 2828 39506 2884 40236
rect 2940 39844 2996 41244
rect 2940 39778 2996 39788
rect 3052 39620 3108 39630
rect 3052 39526 3108 39564
rect 2828 39454 2830 39506
rect 2882 39454 2884 39506
rect 2828 39442 2884 39454
rect 2604 38834 2660 39004
rect 2604 38782 2606 38834
rect 2658 38782 2660 38834
rect 2604 38770 2660 38782
rect 2940 39394 2996 39406
rect 2940 39342 2942 39394
rect 2994 39342 2996 39394
rect 2492 38612 2660 38668
rect 2492 38052 2548 38062
rect 2380 38050 2548 38052
rect 2380 37998 2494 38050
rect 2546 37998 2548 38050
rect 2380 37996 2548 37998
rect 2380 37716 2436 37726
rect 2268 35812 2324 35822
rect 2156 35810 2324 35812
rect 2156 35758 2270 35810
rect 2322 35758 2324 35810
rect 2156 35756 2324 35758
rect 2268 35746 2324 35756
rect 2044 35186 2100 35196
rect 2380 35028 2436 37660
rect 2492 37378 2548 37996
rect 2604 37938 2660 38612
rect 2604 37886 2606 37938
rect 2658 37886 2660 37938
rect 2604 37874 2660 37886
rect 2828 37828 2884 37838
rect 2828 37734 2884 37772
rect 2604 37492 2660 37502
rect 2604 37398 2660 37436
rect 2492 37326 2494 37378
rect 2546 37326 2548 37378
rect 2492 36482 2548 37326
rect 2604 37044 2660 37054
rect 2604 36950 2660 36988
rect 2492 36430 2494 36482
rect 2546 36430 2548 36482
rect 2492 35922 2548 36430
rect 2716 36482 2772 36494
rect 2716 36430 2718 36482
rect 2770 36430 2772 36482
rect 2716 36036 2772 36430
rect 2940 36372 2996 39342
rect 2940 36306 2996 36316
rect 3052 38052 3108 38062
rect 3164 38052 3220 41916
rect 3052 38050 3220 38052
rect 3052 37998 3054 38050
rect 3106 37998 3220 38050
rect 3052 37996 3220 37998
rect 2716 35970 2772 35980
rect 2940 36036 2996 36046
rect 2492 35870 2494 35922
rect 2546 35870 2548 35922
rect 2492 35858 2548 35870
rect 2604 35924 2660 35934
rect 2604 35830 2660 35868
rect 2828 35924 2884 35934
rect 2940 35924 2996 35980
rect 2828 35922 2996 35924
rect 2828 35870 2830 35922
rect 2882 35870 2996 35922
rect 2828 35868 2996 35870
rect 2716 35700 2772 35710
rect 2716 35606 2772 35644
rect 2828 35476 2884 35868
rect 2380 34962 2436 34972
rect 2492 35420 2884 35476
rect 2940 35700 2996 35710
rect 2044 34804 2100 34814
rect 2268 34804 2324 34814
rect 2492 34804 2548 35420
rect 2716 35252 2772 35262
rect 2716 34914 2772 35196
rect 2828 35028 2884 35038
rect 2940 35028 2996 35644
rect 3052 35588 3108 37996
rect 3164 37156 3220 37166
rect 3164 37062 3220 37100
rect 3276 37044 3332 42700
rect 3500 42194 3556 43598
rect 3612 43652 3668 47182
rect 3724 47124 3780 47134
rect 3724 46786 3780 47068
rect 3724 46734 3726 46786
rect 3778 46734 3780 46786
rect 3724 46722 3780 46734
rect 3948 46676 4004 47404
rect 4060 47124 4116 48078
rect 6076 48132 6132 48142
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4060 47058 4116 47068
rect 4508 47346 4564 47358
rect 4508 47294 4510 47346
rect 4562 47294 4564 47346
rect 4508 46900 4564 47294
rect 4508 46834 4564 46844
rect 4844 46788 4900 46798
rect 4844 46694 4900 46732
rect 4508 46676 4564 46686
rect 3948 46674 4564 46676
rect 3948 46622 3950 46674
rect 4002 46622 4510 46674
rect 4562 46622 4564 46674
rect 3948 46620 4564 46622
rect 3836 46562 3892 46574
rect 3836 46510 3838 46562
rect 3890 46510 3892 46562
rect 3836 45556 3892 46510
rect 3948 45890 4004 46620
rect 4508 46610 4564 46620
rect 5964 46562 6020 46574
rect 5964 46510 5966 46562
rect 6018 46510 6020 46562
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 3948 45838 3950 45890
rect 4002 45838 4004 45890
rect 3948 45826 4004 45838
rect 4508 45780 4564 45790
rect 4508 45686 4564 45724
rect 3836 45500 4228 45556
rect 4172 45444 4228 45500
rect 4172 45106 4228 45388
rect 4172 45054 4174 45106
rect 4226 45054 4228 45106
rect 4172 45042 4228 45054
rect 3724 44996 3780 45006
rect 3780 44940 4004 44996
rect 3724 44902 3780 44940
rect 3612 43586 3668 43596
rect 3500 42142 3502 42194
rect 3554 42142 3556 42194
rect 3500 42130 3556 42142
rect 3388 40402 3444 40414
rect 3388 40350 3390 40402
rect 3442 40350 3444 40402
rect 3388 40292 3444 40350
rect 3388 40226 3444 40236
rect 3948 39618 4004 44940
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5740 44212 5796 44222
rect 5404 44210 5796 44212
rect 5404 44158 5742 44210
rect 5794 44158 5796 44210
rect 5404 44156 5796 44158
rect 4844 43652 4900 43662
rect 4844 43538 4900 43596
rect 5292 43652 5348 43662
rect 5292 43558 5348 43596
rect 4844 43486 4846 43538
rect 4898 43486 4900 43538
rect 4844 43474 4900 43486
rect 4060 43426 4116 43438
rect 4396 43428 4452 43438
rect 4060 43374 4062 43426
rect 4114 43374 4116 43426
rect 4060 42196 4116 43374
rect 4060 42130 4116 42140
rect 4284 43426 4452 43428
rect 4284 43374 4398 43426
rect 4450 43374 4452 43426
rect 4284 43372 4452 43374
rect 4060 41860 4116 41870
rect 4060 41766 4116 41804
rect 4284 40292 4340 43372
rect 4396 43362 4452 43372
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 5292 41972 5348 41982
rect 5404 41972 5460 44156
rect 5740 44146 5796 44156
rect 5852 43428 5908 43438
rect 5852 43334 5908 43372
rect 5292 41970 5796 41972
rect 5292 41918 5294 41970
rect 5346 41918 5796 41970
rect 5292 41916 5796 41918
rect 5292 41906 5348 41916
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5740 41188 5796 41916
rect 5852 41188 5908 41198
rect 5740 41186 5908 41188
rect 5740 41134 5854 41186
rect 5906 41134 5908 41186
rect 5740 41132 5908 41134
rect 4732 40516 4788 40526
rect 5180 40516 5236 40526
rect 4732 40514 4900 40516
rect 4732 40462 4734 40514
rect 4786 40462 4900 40514
rect 4732 40460 4900 40462
rect 4732 40450 4788 40460
rect 4284 40226 4340 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4844 39956 4900 40460
rect 5068 40404 5124 40414
rect 4956 39956 5012 39966
rect 4844 39900 4956 39956
rect 3948 39566 3950 39618
rect 4002 39566 4004 39618
rect 3388 39508 3444 39518
rect 3388 38948 3444 39452
rect 3500 39396 3556 39406
rect 3500 39302 3556 39340
rect 3836 39172 3892 39182
rect 3612 39060 3668 39070
rect 3500 38948 3556 38958
rect 3388 38892 3500 38948
rect 3500 38854 3556 38892
rect 3612 37828 3668 39004
rect 3836 39058 3892 39116
rect 3836 39006 3838 39058
rect 3890 39006 3892 39058
rect 3836 38994 3892 39006
rect 3948 38836 4004 39566
rect 3948 38770 4004 38780
rect 4172 39844 4228 39854
rect 4060 38612 4116 38622
rect 4060 38050 4116 38556
rect 4060 37998 4062 38050
rect 4114 37998 4116 38050
rect 4060 37986 4116 37998
rect 4172 38050 4228 39788
rect 4844 39508 4900 39900
rect 4956 39890 5012 39900
rect 5068 39618 5124 40348
rect 5068 39566 5070 39618
rect 5122 39566 5124 39618
rect 5068 39554 5124 39566
rect 4284 39452 4900 39508
rect 4956 39506 5012 39518
rect 4956 39454 4958 39506
rect 5010 39454 5012 39506
rect 4284 39172 4340 39452
rect 4956 39396 5012 39454
rect 5180 39396 5236 40460
rect 5292 40402 5348 40414
rect 5292 40350 5294 40402
rect 5346 40350 5348 40402
rect 5292 40292 5348 40350
rect 5740 40404 5796 41132
rect 5852 41122 5908 41132
rect 5740 40310 5796 40348
rect 5292 40226 5348 40236
rect 5404 40290 5460 40302
rect 5404 40238 5406 40290
rect 5458 40238 5460 40290
rect 4956 39340 5236 39396
rect 4284 39058 4340 39116
rect 4284 39006 4286 39058
rect 4338 39006 4340 39058
rect 4284 38994 4340 39006
rect 4956 39172 5012 39182
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4956 38274 5012 39116
rect 5180 38836 5236 38846
rect 5180 38742 5236 38780
rect 5404 38668 5460 40238
rect 5628 39508 5684 39518
rect 5628 38948 5684 39452
rect 5740 39060 5796 39070
rect 5740 38966 5796 39004
rect 5628 38854 5684 38892
rect 5964 38668 6020 46510
rect 6076 40516 6132 48076
rect 6412 47908 6468 49646
rect 6972 49698 7028 49710
rect 6972 49646 6974 49698
rect 7026 49646 7028 49698
rect 6412 47842 6468 47852
rect 6636 49138 6692 49150
rect 6636 49086 6638 49138
rect 6690 49086 6692 49138
rect 6636 48244 6692 49086
rect 6636 47458 6692 48188
rect 6636 47406 6638 47458
rect 6690 47406 6692 47458
rect 6188 47346 6244 47358
rect 6188 47294 6190 47346
rect 6242 47294 6244 47346
rect 6188 45556 6244 47294
rect 6412 46788 6468 46798
rect 6636 46788 6692 47406
rect 6412 46786 6692 46788
rect 6412 46734 6414 46786
rect 6466 46734 6692 46786
rect 6412 46732 6692 46734
rect 6412 46722 6468 46732
rect 6972 46676 7028 49646
rect 7084 49026 7140 50652
rect 7196 50764 7308 50820
rect 7196 49924 7252 50764
rect 7308 50726 7364 50764
rect 7644 50370 7700 50382
rect 7644 50318 7646 50370
rect 7698 50318 7700 50370
rect 7532 49924 7588 49934
rect 7196 49922 7588 49924
rect 7196 49870 7198 49922
rect 7250 49870 7534 49922
rect 7586 49870 7588 49922
rect 7196 49868 7588 49870
rect 7196 49858 7252 49868
rect 7532 49858 7588 49868
rect 7084 48974 7086 49026
rect 7138 48974 7140 49026
rect 7084 48962 7140 48974
rect 7084 48354 7140 48366
rect 7084 48302 7086 48354
rect 7138 48302 7140 48354
rect 7084 48244 7140 48302
rect 7084 48178 7140 48188
rect 7196 48242 7252 48254
rect 7196 48190 7198 48242
rect 7250 48190 7252 48242
rect 7196 48132 7252 48190
rect 7196 48076 7476 48132
rect 6748 46674 7028 46676
rect 6748 46622 6974 46674
rect 7026 46622 7028 46674
rect 6748 46620 7028 46622
rect 6188 45490 6244 45500
rect 6524 45778 6580 45790
rect 6524 45726 6526 45778
rect 6578 45726 6580 45778
rect 6524 45444 6580 45726
rect 6524 45378 6580 45388
rect 6636 45666 6692 45678
rect 6636 45614 6638 45666
rect 6690 45614 6692 45666
rect 6524 44772 6580 44782
rect 6412 44716 6524 44772
rect 6188 43652 6244 43662
rect 6188 43558 6244 43596
rect 6412 43650 6468 44716
rect 6524 44706 6580 44716
rect 6636 44548 6692 45614
rect 6748 45668 6804 46620
rect 6972 46610 7028 46620
rect 7084 48018 7140 48030
rect 7084 47966 7086 48018
rect 7138 47966 7140 48018
rect 6860 45892 6916 45902
rect 7084 45892 7140 47966
rect 7420 47460 7476 48076
rect 7532 47460 7588 47470
rect 7420 47404 7532 47460
rect 7532 47394 7588 47404
rect 7308 47348 7364 47358
rect 7308 47346 7476 47348
rect 7308 47294 7310 47346
rect 7362 47294 7476 47346
rect 7308 47292 7476 47294
rect 7308 47282 7364 47292
rect 7308 47124 7364 47134
rect 7308 46674 7364 47068
rect 7308 46622 7310 46674
rect 7362 46622 7364 46674
rect 7308 46610 7364 46622
rect 7420 46676 7476 47292
rect 7476 46620 7588 46676
rect 7420 46610 7476 46620
rect 7420 46116 7476 46126
rect 7308 46060 7420 46116
rect 6860 45890 7140 45892
rect 6860 45838 6862 45890
rect 6914 45838 7140 45890
rect 6860 45836 7140 45838
rect 6860 45826 6916 45836
rect 7084 45668 7140 45836
rect 6748 45612 6916 45668
rect 6748 45444 6804 45454
rect 6748 44994 6804 45388
rect 6748 44942 6750 44994
rect 6802 44942 6804 44994
rect 6748 44930 6804 44942
rect 6860 45106 6916 45612
rect 7084 45602 7140 45612
rect 7196 45890 7252 45902
rect 7196 45838 7198 45890
rect 7250 45838 7252 45890
rect 6860 45054 6862 45106
rect 6914 45054 6916 45106
rect 6412 43598 6414 43650
rect 6466 43598 6468 43650
rect 6412 43586 6468 43598
rect 6524 44492 6692 44548
rect 6300 43426 6356 43438
rect 6300 43374 6302 43426
rect 6354 43374 6356 43426
rect 6300 42308 6356 43374
rect 6300 42242 6356 42252
rect 6412 42084 6468 42094
rect 6412 41990 6468 42028
rect 6188 40516 6244 40526
rect 6076 40460 6188 40516
rect 6188 40422 6244 40460
rect 6188 40292 6244 40302
rect 6076 39956 6132 39966
rect 6076 39730 6132 39900
rect 6076 39678 6078 39730
rect 6130 39678 6132 39730
rect 6076 39666 6132 39678
rect 6188 38834 6244 40236
rect 6524 39284 6580 44492
rect 6860 44322 6916 45054
rect 6860 44270 6862 44322
rect 6914 44270 6916 44322
rect 6860 44212 6916 44270
rect 6860 44146 6916 44156
rect 6972 45556 7028 45566
rect 6972 45106 7028 45500
rect 6972 45054 6974 45106
rect 7026 45054 7028 45106
rect 6972 43538 7028 45054
rect 7196 44772 7252 45838
rect 7196 44706 7252 44716
rect 6972 43486 6974 43538
rect 7026 43486 7028 43538
rect 6860 43428 6916 43438
rect 6188 38782 6190 38834
rect 6242 38782 6244 38834
rect 6188 38770 6244 38782
rect 6300 39228 6580 39284
rect 6636 43204 6692 43214
rect 6300 38668 6356 39228
rect 6524 38836 6580 38874
rect 6524 38770 6580 38780
rect 5404 38612 5572 38668
rect 5292 38388 5348 38398
rect 4956 38222 4958 38274
rect 5010 38222 5012 38274
rect 4956 38210 5012 38222
rect 5180 38332 5292 38388
rect 4172 37998 4174 38050
rect 4226 37998 4228 38050
rect 4172 37986 4228 37998
rect 4732 38052 4788 38062
rect 4732 37958 4788 37996
rect 4284 37938 4340 37950
rect 4284 37886 4286 37938
rect 4338 37886 4340 37938
rect 3612 37826 4004 37828
rect 3612 37774 3614 37826
rect 3666 37774 4004 37826
rect 3612 37772 4004 37774
rect 3612 37762 3668 37772
rect 3612 37268 3668 37278
rect 3276 36988 3556 37044
rect 3276 36482 3332 36494
rect 3276 36430 3278 36482
rect 3330 36430 3332 36482
rect 3276 36036 3332 36430
rect 3276 35970 3332 35980
rect 3500 35922 3556 36988
rect 3612 36594 3668 37212
rect 3612 36542 3614 36594
rect 3666 36542 3668 36594
rect 3612 36530 3668 36542
rect 3836 36372 3892 36382
rect 3836 36278 3892 36316
rect 3500 35870 3502 35922
rect 3554 35870 3556 35922
rect 3500 35858 3556 35870
rect 3724 35810 3780 35822
rect 3724 35758 3726 35810
rect 3778 35758 3780 35810
rect 3276 35700 3332 35710
rect 3276 35606 3332 35644
rect 3052 35532 3220 35588
rect 2828 35026 2996 35028
rect 2828 34974 2830 35026
rect 2882 34974 2996 35026
rect 2828 34972 2996 34974
rect 3052 35364 3108 35374
rect 2828 34962 2884 34972
rect 2716 34862 2718 34914
rect 2770 34862 2772 34914
rect 2716 34850 2772 34862
rect 2100 34802 2324 34804
rect 2100 34750 2270 34802
rect 2322 34750 2324 34802
rect 2100 34748 2324 34750
rect 2044 34738 2100 34748
rect 2268 34738 2324 34748
rect 2380 34802 2548 34804
rect 2380 34750 2494 34802
rect 2546 34750 2548 34802
rect 2380 34748 2548 34750
rect 2044 34244 2100 34254
rect 2380 34244 2436 34748
rect 2492 34738 2548 34748
rect 2828 34804 2884 34814
rect 2828 34802 2996 34804
rect 2828 34750 2830 34802
rect 2882 34750 2996 34802
rect 2828 34748 2996 34750
rect 2828 34738 2884 34748
rect 2940 34692 2996 34748
rect 2940 34626 2996 34636
rect 2492 34580 2548 34590
rect 2548 34524 2660 34580
rect 2492 34514 2548 34524
rect 2492 34356 2548 34366
rect 2492 34262 2548 34300
rect 2044 34150 2100 34188
rect 2268 34188 2436 34244
rect 2044 33124 2100 33134
rect 2044 33030 2100 33068
rect 2268 31892 2324 34188
rect 2492 33236 2548 33246
rect 2492 33142 2548 33180
rect 2604 33012 2660 34524
rect 3052 33572 3108 35308
rect 3164 34692 3220 35532
rect 3164 34626 3220 34636
rect 3276 35308 3332 35318
rect 3052 33506 3108 33516
rect 3276 33346 3332 35252
rect 3276 33294 3278 33346
rect 3330 33294 3332 33346
rect 3276 33282 3332 33294
rect 3500 34018 3556 34030
rect 3500 33966 3502 34018
rect 3554 33966 3556 34018
rect 2492 32956 2660 33012
rect 2828 33234 2884 33246
rect 2828 33182 2830 33234
rect 2882 33182 2884 33234
rect 2268 31218 2324 31836
rect 2268 31166 2270 31218
rect 2322 31166 2324 31218
rect 2268 31154 2324 31166
rect 2380 32562 2436 32574
rect 2380 32510 2382 32562
rect 2434 32510 2436 32562
rect 2156 30996 2212 31006
rect 2156 30902 2212 30940
rect 2044 30324 2100 30334
rect 2380 30324 2436 32510
rect 2492 31668 2548 32956
rect 2828 32788 2884 33182
rect 3500 33236 3556 33966
rect 3724 33460 3780 35758
rect 3836 35476 3892 35486
rect 3836 35382 3892 35420
rect 3948 34354 4004 37772
rect 4284 36484 4340 37886
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4172 36428 4340 36484
rect 4620 36484 4676 36494
rect 3948 34302 3950 34354
rect 4002 34302 4004 34354
rect 3948 34290 4004 34302
rect 4060 35700 4116 35710
rect 3724 33394 3780 33404
rect 4060 33346 4116 35644
rect 4060 33294 4062 33346
rect 4114 33294 4116 33346
rect 4060 33282 4116 33294
rect 3724 33236 3780 33246
rect 3500 33234 3780 33236
rect 3500 33182 3726 33234
rect 3778 33182 3780 33234
rect 3500 33180 3780 33182
rect 2828 32722 2884 32732
rect 3276 32564 3332 32574
rect 3612 32564 3668 32574
rect 2940 32562 3332 32564
rect 2940 32510 3278 32562
rect 3330 32510 3332 32562
rect 2940 32508 3332 32510
rect 2604 31890 2660 31902
rect 2940 31892 2996 32508
rect 3276 32498 3332 32508
rect 3388 32508 3612 32564
rect 3388 31948 3444 32508
rect 3612 32470 3668 32508
rect 2604 31838 2606 31890
rect 2658 31838 2660 31890
rect 2604 31780 2660 31838
rect 2828 31836 2996 31892
rect 3276 31892 3444 31948
rect 3500 31892 3556 31902
rect 2828 31780 2884 31836
rect 2604 31724 2884 31780
rect 2492 31612 2660 31668
rect 2380 30268 2548 30324
rect 2044 30098 2100 30268
rect 2044 30046 2046 30098
rect 2098 30046 2100 30098
rect 2044 30034 2100 30046
rect 2380 30098 2436 30110
rect 2380 30046 2382 30098
rect 2434 30046 2436 30098
rect 2380 29988 2436 30046
rect 2268 29426 2324 29438
rect 2268 29374 2270 29426
rect 2322 29374 2324 29426
rect 2268 28868 2324 29374
rect 2380 28980 2436 29932
rect 2380 28914 2436 28924
rect 2268 28802 2324 28812
rect 2492 28756 2548 30268
rect 2380 28700 2548 28756
rect 2604 28754 2660 31612
rect 2604 28702 2606 28754
rect 2658 28702 2660 28754
rect 2268 28644 2324 28682
rect 2268 28578 2324 28588
rect 2044 28532 2100 28542
rect 2044 28082 2100 28476
rect 2044 28030 2046 28082
rect 2098 28030 2100 28082
rect 2044 28018 2100 28030
rect 2268 28420 2324 28430
rect 2156 27300 2212 27310
rect 2044 25396 2100 25406
rect 1932 25394 2100 25396
rect 1932 25342 2046 25394
rect 2098 25342 2100 25394
rect 1932 25340 2100 25342
rect 1708 25302 1764 25340
rect 2044 25330 2100 25340
rect 1708 23826 1764 23838
rect 1708 23774 1710 23826
rect 1762 23774 1764 23826
rect 1708 23604 1764 23774
rect 2044 23828 2100 23838
rect 2044 23734 2100 23772
rect 1708 23538 1764 23548
rect 1820 23492 1876 23502
rect 1708 22258 1764 22270
rect 1708 22206 1710 22258
rect 1762 22206 1764 22258
rect 1708 21812 1764 22206
rect 1708 21746 1764 21756
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20020 1764 20526
rect 1820 20188 1876 23436
rect 2044 22260 2100 22270
rect 2156 22260 2212 27244
rect 2044 22258 2212 22260
rect 2044 22206 2046 22258
rect 2098 22206 2212 22258
rect 2044 22204 2212 22206
rect 2044 22194 2100 22204
rect 2268 22148 2324 28364
rect 2156 22092 2324 22148
rect 2156 22036 2212 22092
rect 1932 21980 2212 22036
rect 1932 20468 1988 21980
rect 2380 21812 2436 28700
rect 2604 28690 2660 28702
rect 2716 29986 2772 29998
rect 2716 29934 2718 29986
rect 2770 29934 2772 29986
rect 2716 28644 2772 29934
rect 2828 29540 2884 31724
rect 3052 31780 3108 31790
rect 3052 31686 3108 31724
rect 3052 31108 3108 31118
rect 3052 31014 3108 31052
rect 3164 29988 3220 29998
rect 3164 29894 3220 29932
rect 3276 29540 3332 31892
rect 3500 31798 3556 31836
rect 3388 31108 3444 31118
rect 3388 30882 3444 31052
rect 3500 30996 3556 31006
rect 3724 30996 3780 33180
rect 3836 33124 3892 33134
rect 3836 33030 3892 33068
rect 4172 33012 4228 36428
rect 4284 36260 4340 36270
rect 4284 36166 4340 36204
rect 4620 35922 4676 36428
rect 4844 36260 4900 36270
rect 4844 36166 4900 36204
rect 4620 35870 4622 35922
rect 4674 35870 4676 35922
rect 4620 35858 4676 35870
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4396 34356 4452 34366
rect 4284 34300 4396 34356
rect 4284 33346 4340 34300
rect 4396 34290 4452 34300
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4284 33294 4286 33346
rect 4338 33294 4340 33346
rect 4284 33282 4340 33294
rect 4620 33572 4676 33582
rect 4620 33346 4676 33516
rect 4620 33294 4622 33346
rect 4674 33294 4676 33346
rect 4620 33282 4676 33294
rect 5068 33348 5124 33358
rect 5068 33254 5124 33292
rect 3948 32956 4228 33012
rect 4508 33234 4564 33246
rect 4508 33182 4510 33234
rect 4562 33182 4564 33234
rect 3948 32900 4004 32956
rect 3500 30994 3780 30996
rect 3500 30942 3502 30994
rect 3554 30942 3780 30994
rect 3500 30940 3780 30942
rect 3500 30930 3556 30940
rect 3388 30830 3390 30882
rect 3442 30830 3444 30882
rect 3388 30818 3444 30830
rect 3724 30212 3780 30940
rect 3724 30146 3780 30156
rect 3836 32844 4004 32900
rect 2828 29538 2996 29540
rect 2828 29486 2830 29538
rect 2882 29486 2996 29538
rect 2828 29484 2996 29486
rect 2828 29474 2884 29484
rect 2828 28644 2884 28654
rect 2716 28642 2884 28644
rect 2716 28590 2830 28642
rect 2882 28590 2884 28642
rect 2716 28588 2884 28590
rect 2828 28578 2884 28588
rect 2492 28532 2548 28542
rect 2492 28530 2660 28532
rect 2492 28478 2494 28530
rect 2546 28478 2660 28530
rect 2492 28476 2660 28478
rect 2492 28466 2548 28476
rect 2492 27748 2548 27758
rect 2492 27654 2548 27692
rect 2492 25396 2548 25406
rect 2492 25302 2548 25340
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 2044 21756 2436 21812
rect 2492 22146 2548 22158
rect 2492 22094 2494 22146
rect 2546 22094 2548 22146
rect 2492 21812 2548 22094
rect 2044 20690 2100 21756
rect 2492 21746 2548 21756
rect 2604 21140 2660 28476
rect 2716 28420 2772 28430
rect 2940 28420 2996 29484
rect 3276 29474 3332 29484
rect 3388 29540 3444 29550
rect 3388 28644 3444 29484
rect 3836 28754 3892 32844
rect 4508 32340 4564 33182
rect 5180 32786 5236 38332
rect 5292 38322 5348 38332
rect 5404 35028 5460 35038
rect 5180 32734 5182 32786
rect 5234 32734 5236 32786
rect 5180 32722 5236 32734
rect 5292 34692 5348 34702
rect 5292 32676 5348 34636
rect 5404 34356 5460 34972
rect 5404 34262 5460 34300
rect 5404 32676 5460 32686
rect 5292 32674 5460 32676
rect 5292 32622 5406 32674
rect 5458 32622 5460 32674
rect 5292 32620 5460 32622
rect 5404 32610 5460 32620
rect 4956 32564 5012 32574
rect 4956 32470 5012 32508
rect 4284 32284 4564 32340
rect 3948 31556 4004 31566
rect 3948 31462 4004 31500
rect 4284 30994 4340 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5516 31556 5572 38612
rect 5740 38612 6020 38668
rect 6188 38612 6356 38668
rect 6412 38724 6468 38734
rect 6412 38612 6580 38668
rect 5628 38050 5684 38062
rect 5628 37998 5630 38050
rect 5682 37998 5684 38050
rect 5628 37828 5684 37998
rect 5628 37762 5684 37772
rect 5740 36482 5796 38612
rect 6188 37826 6244 38612
rect 6188 37774 6190 37826
rect 6242 37774 6244 37826
rect 6188 37156 6244 37774
rect 6524 38050 6580 38612
rect 6524 37998 6526 38050
rect 6578 37998 6580 38050
rect 6300 37492 6356 37502
rect 6524 37492 6580 37998
rect 6300 37490 6580 37492
rect 6300 37438 6302 37490
rect 6354 37438 6580 37490
rect 6300 37436 6580 37438
rect 6300 37426 6356 37436
rect 6188 37100 6468 37156
rect 5740 36430 5742 36482
rect 5794 36430 5796 36482
rect 5740 35922 5796 36430
rect 5964 36372 6020 36382
rect 6020 36316 6132 36372
rect 5964 36278 6020 36316
rect 5740 35870 5742 35922
rect 5794 35870 5796 35922
rect 5740 35858 5796 35870
rect 5628 34802 5684 34814
rect 5628 34750 5630 34802
rect 5682 34750 5684 34802
rect 5628 32004 5684 34750
rect 5628 31938 5684 31948
rect 5852 34018 5908 34030
rect 5852 33966 5854 34018
rect 5906 33966 5908 34018
rect 5852 31892 5908 33966
rect 5964 33348 6020 33358
rect 5964 33254 6020 33292
rect 5964 31892 6020 31902
rect 5852 31836 5964 31892
rect 5964 31826 6020 31836
rect 6076 31668 6132 36316
rect 6300 35586 6356 35598
rect 6300 35534 6302 35586
rect 6354 35534 6356 35586
rect 6300 35140 6356 35534
rect 6300 35074 6356 35084
rect 6188 34916 6244 34926
rect 6412 34916 6468 37100
rect 6524 34916 6580 34926
rect 6412 34914 6580 34916
rect 6412 34862 6526 34914
rect 6578 34862 6580 34914
rect 6412 34860 6580 34862
rect 6188 34822 6244 34860
rect 6524 34850 6580 34860
rect 6412 34244 6468 34254
rect 6636 34244 6692 43148
rect 6860 41076 6916 43372
rect 6972 42084 7028 43486
rect 6972 42018 7028 42028
rect 7084 42754 7140 42766
rect 7084 42702 7086 42754
rect 7138 42702 7140 42754
rect 6860 41074 7028 41076
rect 6860 41022 6862 41074
rect 6914 41022 7028 41074
rect 6860 41020 7028 41022
rect 6860 41010 6916 41020
rect 6972 40516 7028 41020
rect 6972 37938 7028 40460
rect 7084 38948 7140 42702
rect 7308 42420 7364 46060
rect 7420 46050 7476 46060
rect 7420 43652 7476 43662
rect 7420 43558 7476 43596
rect 7308 42364 7476 42420
rect 7308 42196 7364 42206
rect 7308 41970 7364 42140
rect 7308 41918 7310 41970
rect 7362 41918 7364 41970
rect 7308 41906 7364 41918
rect 7308 40964 7364 40974
rect 7084 38854 7140 38892
rect 7196 40962 7364 40964
rect 7196 40910 7310 40962
rect 7362 40910 7364 40962
rect 7196 40908 7364 40910
rect 6972 37886 6974 37938
rect 7026 37886 7028 37938
rect 6972 37874 7028 37886
rect 6860 37826 6916 37838
rect 6860 37774 6862 37826
rect 6914 37774 6916 37826
rect 6748 36372 6804 36382
rect 6748 36278 6804 36316
rect 6412 32564 6468 34188
rect 6524 34188 6692 34244
rect 6748 35252 6804 35262
rect 6524 33796 6580 34188
rect 6636 34020 6692 34030
rect 6748 34020 6804 35196
rect 6636 34018 6804 34020
rect 6636 33966 6638 34018
rect 6690 33966 6804 34018
rect 6636 33964 6804 33966
rect 6636 33954 6692 33964
rect 6524 33740 6692 33796
rect 6524 32564 6580 32574
rect 6412 32562 6580 32564
rect 6412 32510 6526 32562
rect 6578 32510 6580 32562
rect 6412 32508 6580 32510
rect 6524 32498 6580 32508
rect 5516 31490 5572 31500
rect 5964 31612 6132 31668
rect 6524 32340 6580 32350
rect 4396 31108 4452 31118
rect 4396 31014 4452 31052
rect 5628 31108 5684 31118
rect 5628 31106 5796 31108
rect 5628 31054 5630 31106
rect 5682 31054 5796 31106
rect 5628 31052 5796 31054
rect 5628 31042 5684 31052
rect 4284 30942 4286 30994
rect 4338 30942 4340 30994
rect 4284 30436 4340 30942
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30380 4788 30436
rect 4732 30210 4788 30380
rect 4732 30158 4734 30210
rect 4786 30158 4788 30210
rect 4732 30146 4788 30158
rect 4172 30100 4228 30110
rect 4172 30006 4228 30044
rect 5068 30100 5124 30110
rect 5068 30006 5124 30044
rect 4620 29988 4676 29998
rect 4956 29988 5012 29998
rect 4620 29986 5012 29988
rect 4620 29934 4622 29986
rect 4674 29934 4958 29986
rect 5010 29934 5012 29986
rect 4620 29932 5012 29934
rect 4620 29922 4676 29932
rect 4620 29428 4676 29438
rect 4620 29334 4676 29372
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 3836 28702 3838 28754
rect 3890 28702 3892 28754
rect 3836 28690 3892 28702
rect 3388 28578 3444 28588
rect 3948 28644 4004 28654
rect 3948 28550 4004 28588
rect 3276 28532 3332 28542
rect 4956 28532 5012 29932
rect 5740 29876 5796 31052
rect 5852 29988 5908 29998
rect 5852 29894 5908 29932
rect 5740 29810 5796 29820
rect 5964 29764 6020 31612
rect 6076 31332 6132 31342
rect 6076 29988 6132 31276
rect 6300 30882 6356 30894
rect 6300 30830 6302 30882
rect 6354 30830 6356 30882
rect 6188 30324 6244 30334
rect 6188 30210 6244 30268
rect 6188 30158 6190 30210
rect 6242 30158 6244 30210
rect 6188 30146 6244 30158
rect 6076 29932 6244 29988
rect 5852 29708 6020 29764
rect 5740 29426 5796 29438
rect 5740 29374 5742 29426
rect 5794 29374 5796 29426
rect 5740 28644 5796 29374
rect 5740 28578 5796 28588
rect 5180 28532 5236 28542
rect 4956 28476 5124 28532
rect 3276 28438 3332 28476
rect 2716 28418 2940 28420
rect 2716 28366 2718 28418
rect 2770 28366 2940 28418
rect 2716 28364 2940 28366
rect 2716 28354 2772 28364
rect 2940 28326 2996 28364
rect 3500 28420 3556 28430
rect 3500 28326 3556 28364
rect 3724 28418 3780 28430
rect 3724 28366 3726 28418
rect 3778 28366 3780 28418
rect 3724 27636 3780 28366
rect 4732 28308 4788 28318
rect 4732 28082 4788 28252
rect 4732 28030 4734 28082
rect 4786 28030 4788 28082
rect 4732 28018 4788 28030
rect 4172 27972 4228 27982
rect 4172 27878 4228 27916
rect 4956 27972 5012 27982
rect 4956 27878 5012 27916
rect 3724 27580 3892 27636
rect 3724 27300 3780 27310
rect 3724 27186 3780 27244
rect 3724 27134 3726 27186
rect 3778 27134 3780 27186
rect 3724 27122 3780 27134
rect 3500 26962 3556 26974
rect 3500 26910 3502 26962
rect 3554 26910 3556 26962
rect 3500 26852 3556 26910
rect 3500 26786 3556 26796
rect 3724 26852 3780 26862
rect 3724 26758 3780 26796
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 2044 20626 2100 20638
rect 2380 21084 2660 21140
rect 1932 20412 2324 20468
rect 2268 20188 2324 20412
rect 1820 20132 2100 20188
rect 1708 19954 1764 19964
rect 2044 18674 2100 20132
rect 2044 18622 2046 18674
rect 2098 18622 2100 18674
rect 2044 18610 2100 18622
rect 2156 20132 2324 20188
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18228 1764 18398
rect 1708 18162 1764 18172
rect 2044 17108 2100 17118
rect 2156 17108 2212 20132
rect 2044 17106 2212 17108
rect 2044 17054 2046 17106
rect 2098 17054 2212 17106
rect 2044 17052 2212 17054
rect 2044 17042 2100 17052
rect 1708 16882 1764 16894
rect 2380 16884 2436 21084
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 2492 20020 2548 20526
rect 2492 19954 2548 19964
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2492 18228 2548 18286
rect 2492 18162 2548 18172
rect 1708 16830 1710 16882
rect 1762 16830 1764 16882
rect 1708 16436 1764 16830
rect 1708 16370 1764 16380
rect 2044 16828 2436 16884
rect 2492 16882 2548 16894
rect 2492 16830 2494 16882
rect 2546 16830 2548 16882
rect 1820 15764 1876 15774
rect 1876 15708 1988 15764
rect 1820 15698 1876 15708
rect 1708 15314 1764 15326
rect 1708 15262 1710 15314
rect 1762 15262 1764 15314
rect 1708 14644 1764 15262
rect 1708 14578 1764 14588
rect 1708 12852 1764 12862
rect 1708 12758 1764 12796
rect 1708 11282 1764 11294
rect 1708 11230 1710 11282
rect 1762 11230 1764 11282
rect 1708 11060 1764 11230
rect 1932 11284 1988 15708
rect 2044 15538 2100 16828
rect 2492 16436 2548 16830
rect 2492 16370 2548 16380
rect 2044 15486 2046 15538
rect 2098 15486 2100 15538
rect 2044 15474 2100 15486
rect 2492 15202 2548 15214
rect 2492 15150 2494 15202
rect 2546 15150 2548 15202
rect 2492 14644 2548 15150
rect 2492 14578 2548 14588
rect 2044 13412 2100 13422
rect 2044 12850 2100 13356
rect 3836 13412 3892 27580
rect 5068 27524 5124 28476
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 5068 27458 5124 27468
rect 5180 28082 5236 28476
rect 5740 28308 5796 28318
rect 5180 28030 5182 28082
rect 5234 28030 5236 28082
rect 4476 27402 4740 27412
rect 4620 27300 4676 27310
rect 4620 27188 4676 27244
rect 4284 27186 4676 27188
rect 4284 27134 4622 27186
rect 4674 27134 4676 27186
rect 4284 27132 4676 27134
rect 3948 27076 4004 27086
rect 3948 26982 4004 27020
rect 4284 27074 4340 27132
rect 4620 27122 4676 27132
rect 4284 27022 4286 27074
rect 4338 27022 4340 27074
rect 4284 27010 4340 27022
rect 5180 27076 5236 28030
rect 5516 28084 5572 28094
rect 5292 27860 5348 27870
rect 5292 27746 5348 27804
rect 5516 27858 5572 28028
rect 5516 27806 5518 27858
rect 5570 27806 5572 27858
rect 5516 27794 5572 27806
rect 5628 27972 5684 27982
rect 5292 27694 5294 27746
rect 5346 27694 5348 27746
rect 5292 27682 5348 27694
rect 5180 26908 5236 27020
rect 5180 26852 5572 26908
rect 5516 26290 5572 26852
rect 5516 26238 5518 26290
rect 5570 26238 5572 26290
rect 5516 26226 5572 26238
rect 5068 26068 5124 26078
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 3836 13346 3892 13356
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2044 12798 2046 12850
rect 2098 12798 2100 12850
rect 2044 12786 2100 12798
rect 2492 12852 2548 12862
rect 2492 12758 2548 12796
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 2044 11284 2100 11294
rect 1932 11282 2100 11284
rect 1932 11230 2046 11282
rect 2098 11230 2100 11282
rect 1932 11228 2100 11230
rect 2044 11218 2100 11228
rect 1708 10994 1764 11004
rect 2492 11170 2548 11182
rect 2492 11118 2494 11170
rect 2546 11118 2548 11170
rect 2492 11060 2548 11118
rect 2492 10994 2548 11004
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 1708 9714 1764 9726
rect 1708 9662 1710 9714
rect 1762 9662 1764 9714
rect 1708 9268 1764 9662
rect 2044 9716 2100 9726
rect 2044 9622 2100 9660
rect 2492 9602 2548 9614
rect 2492 9550 2494 9602
rect 2546 9550 2548 9602
rect 1708 9202 1764 9212
rect 2044 9492 2100 9502
rect 1708 8146 1764 8158
rect 1708 8094 1710 8146
rect 1762 8094 1764 8146
rect 1708 8036 1764 8094
rect 2044 8146 2100 9436
rect 2492 9268 2548 9550
rect 2492 9202 2548 9212
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 2044 8094 2046 8146
rect 2098 8094 2100 8146
rect 2044 8082 2100 8094
rect 1708 7476 1764 7980
rect 2492 8036 2548 8046
rect 2492 7942 2548 7980
rect 1708 7410 1764 7420
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 2380 6804 2436 6814
rect 1708 5906 1764 5918
rect 1708 5854 1710 5906
rect 1762 5854 1764 5906
rect 1708 5684 1764 5854
rect 2156 5908 2212 5918
rect 2156 5794 2212 5852
rect 2156 5742 2158 5794
rect 2210 5742 2212 5794
rect 2156 5730 2212 5742
rect 1708 5236 1764 5628
rect 1820 5236 1876 5246
rect 1708 5234 1876 5236
rect 1708 5182 1822 5234
rect 1874 5182 1876 5234
rect 1708 5180 1876 5182
rect 1820 5170 1876 5180
rect 2044 4564 2100 4574
rect 1596 4562 2100 4564
rect 1596 4510 2046 4562
rect 2098 4510 2100 4562
rect 1596 4508 2100 4510
rect 2044 4498 2100 4508
rect 1708 4338 1764 4350
rect 1708 4286 1710 4338
rect 1762 4286 1764 4338
rect 1708 3892 1764 4286
rect 1708 3826 1764 3836
rect 2268 3668 2324 3678
rect 2380 3668 2436 6748
rect 5068 6804 5124 26012
rect 5628 9492 5684 27916
rect 5740 27858 5796 28252
rect 5740 27806 5742 27858
rect 5794 27806 5796 27858
rect 5740 27794 5796 27806
rect 5852 27074 5908 29708
rect 6188 29650 6244 29932
rect 6188 29598 6190 29650
rect 6242 29598 6244 29650
rect 6188 29586 6244 29598
rect 6076 29540 6132 29550
rect 6076 28754 6132 29484
rect 6076 28702 6078 28754
rect 6130 28702 6132 28754
rect 5852 27022 5854 27074
rect 5906 27022 5908 27074
rect 5852 26404 5908 27022
rect 5964 27970 6020 27982
rect 5964 27918 5966 27970
rect 6018 27918 6020 27970
rect 5964 26516 6020 27918
rect 5964 26450 6020 26460
rect 5852 26292 5908 26348
rect 5964 26292 6020 26302
rect 5852 26290 6020 26292
rect 5852 26238 5966 26290
rect 6018 26238 6020 26290
rect 5852 26236 6020 26238
rect 5964 26226 6020 26236
rect 5964 26068 6020 26078
rect 6076 26068 6132 28702
rect 6188 29428 6244 29438
rect 6188 26908 6244 29372
rect 6300 28644 6356 30830
rect 6524 30322 6580 32284
rect 6524 30270 6526 30322
rect 6578 30270 6580 30322
rect 6524 30258 6580 30270
rect 6412 30212 6468 30222
rect 6636 30212 6692 33740
rect 6636 30156 6804 30212
rect 6412 30118 6468 30156
rect 6636 29988 6692 29998
rect 6636 29894 6692 29932
rect 6748 29764 6804 30156
rect 6636 29708 6804 29764
rect 6860 30210 6916 37774
rect 7084 37828 7140 37838
rect 7084 36594 7140 37772
rect 7084 36542 7086 36594
rect 7138 36542 7140 36594
rect 7084 36530 7140 36542
rect 7196 36706 7252 40908
rect 7308 40898 7364 40908
rect 7420 40180 7476 42364
rect 7532 42308 7588 46620
rect 7644 45892 7700 50318
rect 7980 49700 8036 49710
rect 7868 47460 7924 47470
rect 7980 47460 8036 49644
rect 8204 48916 8260 55412
rect 10444 53506 10500 55412
rect 12348 55412 12516 55468
rect 13692 55412 14420 55468
rect 16380 55412 16436 55422
rect 11788 55188 11844 55198
rect 11788 55094 11844 55132
rect 11900 55076 11956 55086
rect 11900 55074 12292 55076
rect 11900 55022 11902 55074
rect 11954 55022 12292 55074
rect 11900 55020 12292 55022
rect 11900 55010 11956 55020
rect 12236 54404 12292 55020
rect 12348 54628 12404 55412
rect 13580 55300 13636 55310
rect 13580 55206 13636 55244
rect 12348 54562 12404 54572
rect 12460 54796 13188 54852
rect 12460 54514 12516 54796
rect 12796 54628 12852 54638
rect 12796 54626 12964 54628
rect 12796 54574 12798 54626
rect 12850 54574 12964 54626
rect 12796 54572 12964 54574
rect 12796 54562 12852 54572
rect 12460 54462 12462 54514
rect 12514 54462 12516 54514
rect 12460 54404 12516 54462
rect 12236 54348 12516 54404
rect 12796 53620 12852 53630
rect 10444 53454 10446 53506
rect 10498 53454 10500 53506
rect 9884 53058 9940 53070
rect 9884 53006 9886 53058
rect 9938 53006 9940 53058
rect 8764 52946 8820 52958
rect 8764 52894 8766 52946
rect 8818 52894 8820 52946
rect 8764 52164 8820 52894
rect 9884 52948 9940 53006
rect 8988 52164 9044 52174
rect 8764 52162 9044 52164
rect 8764 52110 8990 52162
rect 9042 52110 9044 52162
rect 8764 52108 9044 52110
rect 9884 52164 9940 52892
rect 10220 52948 10276 52958
rect 10444 52948 10500 53454
rect 10892 53508 10948 53518
rect 10668 53060 10724 53070
rect 10668 52966 10724 53004
rect 10220 52946 10500 52948
rect 10220 52894 10222 52946
rect 10274 52894 10500 52946
rect 10220 52892 10500 52894
rect 10556 52948 10612 52958
rect 10220 52388 10276 52892
rect 10220 52322 10276 52332
rect 10444 52724 10500 52734
rect 10444 52386 10500 52668
rect 10444 52334 10446 52386
rect 10498 52334 10500 52386
rect 10444 52322 10500 52334
rect 10332 52276 10388 52286
rect 9996 52164 10052 52174
rect 9884 52162 10052 52164
rect 9884 52110 9998 52162
rect 10050 52110 10052 52162
rect 9884 52108 10052 52110
rect 8988 51380 9044 52108
rect 9996 52098 10052 52108
rect 10332 52162 10388 52220
rect 10332 52110 10334 52162
rect 10386 52110 10388 52162
rect 10332 52098 10388 52110
rect 10108 51940 10164 51950
rect 10108 51846 10164 51884
rect 10556 51492 10612 52892
rect 10892 52946 10948 53452
rect 11564 53508 11620 53518
rect 11564 53414 11620 53452
rect 12796 53172 12852 53564
rect 12348 53170 12852 53172
rect 12348 53118 12798 53170
rect 12850 53118 12852 53170
rect 12348 53116 12852 53118
rect 12012 53060 12068 53070
rect 11676 53058 12068 53060
rect 11676 53006 12014 53058
rect 12066 53006 12068 53058
rect 11676 53004 12068 53006
rect 10892 52894 10894 52946
rect 10946 52894 10948 52946
rect 10892 52882 10948 52894
rect 11116 52948 11172 52958
rect 11004 52724 11060 52734
rect 10780 52162 10836 52174
rect 10780 52110 10782 52162
rect 10834 52110 10836 52162
rect 10780 51604 10836 52110
rect 10780 51538 10836 51548
rect 10892 51716 10948 51726
rect 10668 51492 10724 51502
rect 10556 51490 10724 51492
rect 10556 51438 10670 51490
rect 10722 51438 10724 51490
rect 10556 51436 10724 51438
rect 10668 51426 10724 51436
rect 10892 51490 10948 51660
rect 10892 51438 10894 51490
rect 10946 51438 10948 51490
rect 10892 51426 10948 51438
rect 11004 51380 11060 52668
rect 11116 52162 11172 52892
rect 11340 52948 11396 52958
rect 11340 52946 11508 52948
rect 11340 52894 11342 52946
rect 11394 52894 11508 52946
rect 11340 52892 11508 52894
rect 11340 52882 11396 52892
rect 11116 52110 11118 52162
rect 11170 52110 11172 52162
rect 11116 52098 11172 52110
rect 11340 52164 11396 52174
rect 11340 52070 11396 52108
rect 11116 51380 11172 51390
rect 11004 51378 11172 51380
rect 11004 51326 11118 51378
rect 11170 51326 11172 51378
rect 11004 51324 11172 51326
rect 8988 51314 9044 51324
rect 11116 51314 11172 51324
rect 11228 51378 11284 51390
rect 11228 51326 11230 51378
rect 11282 51326 11284 51378
rect 10780 51266 10836 51278
rect 10780 51214 10782 51266
rect 10834 51214 10836 51266
rect 10780 49924 10836 51214
rect 11228 50428 11284 51326
rect 11452 50484 11508 52892
rect 11676 52724 11732 53004
rect 12012 52994 12068 53004
rect 12348 53058 12404 53116
rect 12796 53106 12852 53116
rect 12908 53172 12964 54572
rect 13132 54626 13188 54796
rect 13132 54574 13134 54626
rect 13186 54574 13188 54626
rect 13132 54562 13188 54574
rect 13692 54514 13748 55412
rect 16156 55410 16436 55412
rect 16156 55358 16382 55410
rect 16434 55358 16436 55410
rect 16156 55356 16436 55358
rect 14252 55188 14308 55198
rect 14252 55186 14756 55188
rect 14252 55134 14254 55186
rect 14306 55134 14756 55186
rect 14252 55132 14756 55134
rect 14252 55122 14308 55132
rect 14700 54738 14756 55132
rect 15820 54740 15876 54750
rect 14700 54686 14702 54738
rect 14754 54686 14756 54738
rect 14700 54674 14756 54686
rect 15148 54738 15876 54740
rect 15148 54686 15822 54738
rect 15874 54686 15876 54738
rect 15148 54684 15876 54686
rect 15148 54626 15204 54684
rect 15820 54674 15876 54684
rect 15148 54574 15150 54626
rect 15202 54574 15204 54626
rect 15148 54562 15204 54574
rect 13692 54462 13694 54514
rect 13746 54462 13748 54514
rect 13692 54450 13748 54462
rect 14588 54514 14644 54526
rect 14588 54462 14590 54514
rect 14642 54462 14644 54514
rect 13804 54402 13860 54414
rect 13804 54350 13806 54402
rect 13858 54350 13860 54402
rect 13804 53620 13860 54350
rect 13804 53554 13860 53564
rect 12908 53106 12964 53116
rect 12348 53006 12350 53058
rect 12402 53006 12404 53058
rect 12348 52994 12404 53006
rect 11676 52386 11732 52668
rect 12796 52724 12852 52734
rect 11676 52334 11678 52386
rect 11730 52334 11732 52386
rect 11676 52322 11732 52334
rect 12460 52388 12516 52398
rect 11900 52164 11956 52174
rect 12348 52164 12404 52174
rect 11900 52162 12292 52164
rect 11900 52110 11902 52162
rect 11954 52110 12292 52162
rect 11900 52108 12292 52110
rect 11900 52098 11956 52108
rect 11900 51938 11956 51950
rect 11900 51886 11902 51938
rect 11954 51886 11956 51938
rect 11116 50372 11284 50428
rect 11340 50428 11508 50484
rect 11564 51604 11620 51614
rect 11116 50036 11172 50372
rect 11340 50260 11396 50428
rect 11116 49970 11172 49980
rect 11228 50204 11396 50260
rect 10780 49858 10836 49868
rect 8540 49812 8596 49822
rect 8540 49698 8596 49756
rect 8540 49646 8542 49698
rect 8594 49646 8596 49698
rect 8540 49634 8596 49646
rect 8876 49810 8932 49822
rect 8876 49758 8878 49810
rect 8930 49758 8932 49810
rect 8876 49700 8932 49758
rect 10444 49812 10500 49822
rect 11228 49812 11284 50204
rect 11564 50148 11620 51548
rect 11900 51268 11956 51886
rect 12012 51604 12068 51614
rect 12012 51510 12068 51548
rect 11900 51202 11956 51212
rect 12236 50428 12292 52108
rect 12348 52070 12404 52108
rect 11340 50092 11620 50148
rect 11900 50370 11956 50382
rect 12236 50372 12404 50428
rect 11900 50318 11902 50370
rect 11954 50318 11956 50370
rect 11340 50034 11396 50092
rect 11340 49982 11342 50034
rect 11394 49982 11396 50034
rect 11340 49970 11396 49982
rect 11564 49812 11620 49822
rect 11900 49812 11956 50318
rect 12012 50036 12068 50046
rect 12012 49942 12068 49980
rect 12236 49812 12292 49822
rect 11228 49756 11396 49812
rect 10444 49718 10500 49756
rect 8876 49634 8932 49644
rect 10108 49698 10164 49710
rect 10108 49646 10110 49698
rect 10162 49646 10164 49698
rect 8204 48850 8260 48860
rect 9660 48802 9716 48814
rect 9660 48750 9662 48802
rect 9714 48750 9716 48802
rect 8316 48468 8372 48478
rect 7924 47404 8036 47460
rect 8204 47908 8260 47918
rect 7868 47366 7924 47404
rect 7868 46788 7924 46798
rect 7868 46694 7924 46732
rect 8204 46004 8260 47852
rect 8316 47458 8372 48412
rect 9660 48468 9716 48750
rect 10108 48804 10164 49646
rect 11228 49588 11284 49598
rect 10220 49586 11284 49588
rect 10220 49534 11230 49586
rect 11282 49534 11284 49586
rect 10220 49532 11284 49534
rect 10220 49138 10276 49532
rect 10556 49140 10612 49150
rect 10220 49086 10222 49138
rect 10274 49086 10276 49138
rect 10220 49074 10276 49086
rect 10444 49084 10556 49140
rect 10332 48804 10388 48814
rect 10108 48748 10332 48804
rect 10332 48738 10388 48748
rect 9660 48402 9716 48412
rect 9660 48242 9716 48254
rect 9660 48190 9662 48242
rect 9714 48190 9716 48242
rect 8316 47406 8318 47458
rect 8370 47406 8372 47458
rect 8316 47124 8372 47406
rect 8316 47058 8372 47068
rect 8428 47684 8484 47694
rect 8204 45948 8372 46004
rect 7644 45890 8260 45892
rect 7644 45838 7646 45890
rect 7698 45838 8260 45890
rect 7644 45836 8260 45838
rect 7644 45826 7700 45836
rect 8092 45668 8148 45678
rect 8092 45574 8148 45612
rect 7980 45444 8036 45454
rect 7980 45218 8036 45388
rect 8204 45330 8260 45836
rect 8204 45278 8206 45330
rect 8258 45278 8260 45330
rect 8204 45266 8260 45278
rect 7980 45166 7982 45218
rect 8034 45166 8036 45218
rect 7980 45154 8036 45166
rect 7756 45108 7812 45118
rect 7756 45014 7812 45052
rect 8204 44994 8260 45006
rect 8204 44942 8206 44994
rect 8258 44942 8260 44994
rect 8092 44212 8148 44222
rect 8092 44118 8148 44156
rect 7644 43540 7700 43550
rect 7644 42754 7700 43484
rect 7868 43428 7924 43438
rect 7868 43334 7924 43372
rect 7644 42702 7646 42754
rect 7698 42702 7700 42754
rect 7644 42532 7700 42702
rect 7644 42466 7700 42476
rect 7532 42252 8036 42308
rect 7644 42084 7700 42094
rect 7420 39842 7476 40124
rect 7420 39790 7422 39842
rect 7474 39790 7476 39842
rect 7420 39778 7476 39790
rect 7532 41748 7588 41758
rect 7532 39172 7588 41692
rect 7644 41298 7700 42028
rect 7644 41246 7646 41298
rect 7698 41246 7700 41298
rect 7644 41234 7700 41246
rect 7980 39618 8036 42252
rect 7980 39566 7982 39618
rect 8034 39566 8036 39618
rect 7868 39508 7924 39518
rect 7532 39106 7588 39116
rect 7756 39506 7924 39508
rect 7756 39454 7870 39506
rect 7922 39454 7924 39506
rect 7756 39452 7924 39454
rect 7644 38948 7700 38958
rect 7756 38948 7812 39452
rect 7868 39442 7924 39452
rect 7980 39284 8036 39566
rect 7700 38892 7812 38948
rect 7868 39228 8036 39284
rect 8092 41188 8148 41198
rect 7644 38836 7700 38892
rect 7420 38834 7700 38836
rect 7420 38782 7646 38834
rect 7698 38782 7700 38834
rect 7420 38780 7700 38782
rect 7420 38162 7476 38780
rect 7644 38770 7700 38780
rect 7868 38834 7924 39228
rect 7868 38782 7870 38834
rect 7922 38782 7924 38834
rect 7420 38110 7422 38162
rect 7474 38110 7476 38162
rect 7420 38098 7476 38110
rect 7532 38610 7588 38622
rect 7532 38558 7534 38610
rect 7586 38558 7588 38610
rect 7196 36654 7198 36706
rect 7250 36654 7252 36706
rect 7196 35308 7252 36654
rect 7420 37492 7476 37502
rect 7420 37154 7476 37436
rect 7532 37268 7588 38558
rect 7756 38052 7812 38062
rect 7868 38052 7924 38782
rect 7980 38724 8036 38762
rect 7980 38658 8036 38668
rect 7756 38050 7924 38052
rect 7756 37998 7758 38050
rect 7810 37998 7924 38050
rect 7756 37996 7924 37998
rect 7756 37986 7812 37996
rect 7756 37268 7812 37278
rect 7532 37266 7812 37268
rect 7532 37214 7758 37266
rect 7810 37214 7812 37266
rect 7532 37212 7812 37214
rect 7420 37102 7422 37154
rect 7474 37102 7476 37154
rect 7196 35252 7364 35308
rect 7308 34916 7364 35252
rect 7420 35252 7476 37102
rect 7644 35922 7700 37212
rect 7756 37202 7812 37212
rect 7644 35870 7646 35922
rect 7698 35870 7700 35922
rect 7644 35858 7700 35870
rect 7980 36036 8036 36046
rect 7980 35588 8036 35980
rect 8092 35924 8148 41132
rect 8204 39060 8260 44942
rect 8316 43540 8372 45948
rect 8428 44996 8484 47628
rect 8764 47572 8820 47582
rect 8764 47478 8820 47516
rect 9212 47348 9268 47358
rect 9660 47348 9716 48190
rect 9212 47346 9716 47348
rect 9212 47294 9214 47346
rect 9266 47294 9716 47346
rect 9212 47292 9716 47294
rect 10220 48130 10276 48142
rect 10220 48078 10222 48130
rect 10274 48078 10276 48130
rect 9100 46788 9156 46798
rect 9212 46788 9268 47292
rect 10108 47234 10164 47246
rect 10108 47182 10110 47234
rect 10162 47182 10164 47234
rect 9324 46900 9380 46910
rect 9380 46844 9492 46900
rect 9324 46834 9380 46844
rect 9156 46732 9268 46788
rect 9100 46722 9156 46732
rect 8652 45892 8708 45902
rect 8652 45798 8708 45836
rect 9324 45780 9380 45790
rect 9324 45686 9380 45724
rect 8428 44930 8484 44940
rect 8316 43446 8372 43484
rect 8540 44434 8596 44446
rect 8540 44382 8542 44434
rect 8594 44382 8596 44434
rect 8540 43764 8596 44382
rect 8428 42644 8484 42654
rect 8428 42082 8484 42588
rect 8428 42030 8430 42082
rect 8482 42030 8484 42082
rect 8428 42018 8484 42030
rect 8428 40404 8484 40414
rect 8540 40404 8596 43708
rect 8764 43538 8820 43550
rect 8764 43486 8766 43538
rect 8818 43486 8820 43538
rect 8764 43428 8820 43486
rect 9100 43540 9156 43550
rect 9100 43446 9156 43484
rect 8764 43362 8820 43372
rect 8764 42756 8820 42766
rect 8652 42196 8708 42206
rect 8764 42196 8820 42700
rect 8708 42140 8820 42196
rect 8652 42130 8708 42140
rect 8764 41972 8820 42140
rect 8876 42196 8932 42206
rect 8876 42102 8932 42140
rect 8764 41916 9380 41972
rect 8428 40402 8596 40404
rect 8428 40350 8430 40402
rect 8482 40350 8596 40402
rect 8428 40348 8596 40350
rect 8652 41860 8708 41870
rect 8652 40402 8708 41804
rect 9212 41186 9268 41198
rect 9212 41134 9214 41186
rect 9266 41134 9268 41186
rect 9212 40964 9268 41134
rect 9324 41186 9380 41916
rect 9324 41134 9326 41186
rect 9378 41134 9380 41186
rect 9324 41122 9380 41134
rect 9436 40964 9492 46844
rect 9884 46452 9940 46462
rect 9772 46396 9884 46452
rect 9548 45892 9604 45902
rect 9548 41300 9604 45836
rect 9772 45106 9828 46396
rect 9884 46386 9940 46396
rect 9884 46004 9940 46014
rect 9884 45910 9940 45948
rect 9772 45054 9774 45106
rect 9826 45054 9828 45106
rect 9660 44996 9716 45006
rect 9660 41300 9716 44940
rect 9772 44660 9828 45054
rect 9772 44594 9828 44604
rect 9996 45780 10052 45790
rect 9996 43540 10052 45724
rect 10108 44996 10164 47182
rect 10220 47012 10276 48078
rect 10220 45892 10276 46956
rect 10332 46900 10388 46910
rect 10332 46786 10388 46844
rect 10332 46734 10334 46786
rect 10386 46734 10388 46786
rect 10332 46722 10388 46734
rect 10444 46228 10500 49084
rect 10556 49074 10612 49084
rect 10556 48354 10612 48366
rect 10556 48302 10558 48354
rect 10610 48302 10612 48354
rect 10556 47572 10612 48302
rect 10668 48242 10724 48254
rect 10668 48190 10670 48242
rect 10722 48190 10724 48242
rect 10668 48132 10724 48190
rect 10668 48066 10724 48076
rect 10556 47460 10612 47516
rect 10668 47460 10724 47470
rect 10556 47458 10724 47460
rect 10556 47406 10670 47458
rect 10722 47406 10724 47458
rect 10556 47404 10724 47406
rect 10444 46162 10500 46172
rect 10332 45892 10388 45902
rect 10220 45890 10388 45892
rect 10220 45838 10334 45890
rect 10386 45838 10388 45890
rect 10220 45836 10388 45838
rect 10220 45220 10276 45836
rect 10332 45826 10388 45836
rect 10668 45780 10724 47404
rect 10780 46674 10836 49532
rect 11228 49522 11284 49532
rect 11228 49364 11284 49374
rect 11116 48916 11172 48926
rect 11004 48914 11172 48916
rect 11004 48862 11118 48914
rect 11170 48862 11172 48914
rect 11004 48860 11172 48862
rect 11004 48804 11060 48860
rect 11116 48850 11172 48860
rect 11004 47236 11060 48748
rect 11228 48244 11284 49308
rect 11340 49138 11396 49756
rect 11340 49086 11342 49138
rect 11394 49086 11396 49138
rect 11340 49074 11396 49086
rect 11452 49810 12236 49812
rect 11452 49758 11566 49810
rect 11618 49758 12236 49810
rect 11452 49756 12236 49758
rect 11452 49026 11508 49756
rect 11564 49746 11620 49756
rect 11900 49588 11956 49598
rect 11452 48974 11454 49026
rect 11506 48974 11508 49026
rect 11452 48962 11508 48974
rect 11788 49586 11956 49588
rect 11788 49534 11902 49586
rect 11954 49534 11956 49586
rect 11788 49532 11956 49534
rect 11788 48468 11844 49532
rect 11900 49522 11956 49532
rect 11900 49140 11956 49150
rect 12012 49140 12068 49756
rect 12236 49718 12292 49756
rect 11900 49138 12068 49140
rect 11900 49086 11902 49138
rect 11954 49086 12068 49138
rect 11900 49084 12068 49086
rect 11900 49074 11956 49084
rect 11788 48412 11956 48468
rect 11340 48244 11396 48254
rect 11788 48244 11844 48254
rect 11228 48242 11396 48244
rect 11228 48190 11342 48242
rect 11394 48190 11396 48242
rect 11228 48188 11396 48190
rect 11116 47460 11172 47470
rect 11116 47366 11172 47404
rect 11004 47180 11172 47236
rect 11116 47068 11172 47180
rect 10780 46622 10782 46674
rect 10834 46622 10836 46674
rect 10780 46452 10836 46622
rect 10780 46386 10836 46396
rect 10892 47012 11172 47068
rect 10892 46116 10948 47012
rect 10668 45714 10724 45724
rect 10780 46060 10948 46116
rect 10220 45154 10276 45164
rect 10444 45666 10500 45678
rect 10444 45614 10446 45666
rect 10498 45614 10500 45666
rect 10108 44930 10164 44940
rect 10108 44772 10164 44782
rect 10108 44434 10164 44716
rect 10108 44382 10110 44434
rect 10162 44382 10164 44434
rect 10108 44324 10164 44382
rect 10108 44100 10164 44268
rect 10220 44660 10276 44670
rect 10220 44322 10276 44604
rect 10220 44270 10222 44322
rect 10274 44270 10276 44322
rect 10220 44258 10276 44270
rect 10108 44044 10276 44100
rect 9884 43538 10052 43540
rect 9884 43486 9998 43538
rect 10050 43486 10052 43538
rect 9884 43484 10052 43486
rect 9884 42644 9940 43484
rect 9996 43474 10052 43484
rect 10108 43538 10164 43550
rect 10108 43486 10110 43538
rect 10162 43486 10164 43538
rect 10108 42756 10164 43486
rect 10220 43426 10276 44044
rect 10220 43374 10222 43426
rect 10274 43374 10276 43426
rect 10220 43362 10276 43374
rect 10108 42690 10164 42700
rect 9884 42550 9940 42588
rect 10220 42308 10276 42318
rect 9996 41300 10052 41310
rect 9660 41244 9828 41300
rect 9548 41206 9604 41244
rect 8652 40350 8654 40402
rect 8706 40350 8708 40402
rect 8428 40338 8484 40348
rect 8204 38994 8260 39004
rect 8316 39732 8372 39742
rect 8204 38052 8260 38062
rect 8204 37490 8260 37996
rect 8204 37438 8206 37490
rect 8258 37438 8260 37490
rect 8204 37426 8260 37438
rect 8316 36820 8372 39676
rect 8652 39618 8708 40350
rect 8652 39566 8654 39618
rect 8706 39566 8708 39618
rect 8652 39554 8708 39566
rect 8764 40908 9492 40964
rect 9660 41076 9716 41086
rect 9772 41076 9828 41244
rect 9772 41020 9940 41076
rect 9660 40962 9716 41020
rect 9660 40910 9662 40962
rect 9714 40910 9716 40962
rect 8764 40290 8820 40908
rect 9548 40852 9604 40862
rect 8764 40238 8766 40290
rect 8818 40238 8820 40290
rect 8764 39506 8820 40238
rect 8764 39454 8766 39506
rect 8818 39454 8820 39506
rect 8764 39442 8820 39454
rect 9100 40402 9156 40414
rect 9100 40350 9102 40402
rect 9154 40350 9156 40402
rect 8540 38724 8596 38762
rect 8540 38658 8596 38668
rect 8988 37604 9044 37614
rect 8764 37380 8820 37390
rect 8764 37286 8820 37324
rect 8204 36764 8372 36820
rect 8652 37266 8708 37278
rect 8652 37214 8654 37266
rect 8706 37214 8708 37266
rect 8204 36594 8260 36764
rect 8652 36708 8708 37214
rect 8988 37266 9044 37548
rect 8988 37214 8990 37266
rect 9042 37214 9044 37266
rect 8988 37202 9044 37214
rect 8652 36642 8708 36652
rect 8204 36542 8206 36594
rect 8258 36542 8260 36594
rect 8204 36530 8260 36542
rect 8652 36482 8708 36494
rect 8652 36430 8654 36482
rect 8706 36430 8708 36482
rect 8652 36260 8708 36430
rect 8988 36260 9044 36270
rect 8652 36258 9044 36260
rect 8652 36206 8990 36258
rect 9042 36206 9044 36258
rect 8652 36204 9044 36206
rect 8092 35868 8372 35924
rect 8092 35588 8148 35598
rect 7980 35586 8148 35588
rect 7980 35534 8094 35586
rect 8146 35534 8148 35586
rect 7980 35532 8148 35534
rect 8092 35522 8148 35532
rect 7420 35186 7476 35196
rect 8092 34916 8148 34926
rect 7308 34850 7364 34860
rect 7868 34860 8092 34916
rect 7644 34802 7700 34814
rect 7644 34750 7646 34802
rect 7698 34750 7700 34802
rect 7084 34020 7140 34030
rect 7420 34020 7476 34030
rect 7084 34018 7420 34020
rect 7084 33966 7086 34018
rect 7138 33966 7420 34018
rect 7084 33964 7420 33966
rect 7084 33954 7140 33964
rect 7420 33926 7476 33964
rect 7420 33234 7476 33246
rect 7420 33182 7422 33234
rect 7474 33182 7476 33234
rect 7084 33124 7140 33134
rect 7084 32004 7140 33068
rect 7308 32564 7364 32574
rect 7308 32470 7364 32508
rect 6972 31892 7028 31902
rect 6972 30994 7028 31836
rect 6972 30942 6974 30994
rect 7026 30942 7028 30994
rect 6972 30548 7028 30942
rect 6972 30482 7028 30492
rect 6860 30158 6862 30210
rect 6914 30158 6916 30210
rect 6412 29540 6468 29550
rect 6412 29446 6468 29484
rect 6412 28644 6468 28654
rect 6300 28642 6468 28644
rect 6300 28590 6414 28642
rect 6466 28590 6468 28642
rect 6300 28588 6468 28590
rect 6412 28578 6468 28588
rect 6636 28418 6692 29708
rect 6636 28366 6638 28418
rect 6690 28366 6692 28418
rect 6636 28354 6692 28366
rect 6636 27858 6692 27870
rect 6636 27806 6638 27858
rect 6690 27806 6692 27858
rect 6412 27524 6468 27534
rect 6412 27186 6468 27468
rect 6412 27134 6414 27186
rect 6466 27134 6468 27186
rect 6412 27122 6468 27134
rect 6636 27188 6692 27806
rect 6636 27122 6692 27132
rect 6188 26852 6356 26908
rect 6020 26012 6132 26068
rect 5964 26002 6020 26012
rect 6300 21812 6356 26852
rect 6300 21746 6356 21756
rect 6748 26852 6804 26862
rect 6748 9716 6804 26796
rect 6860 26292 6916 30158
rect 7084 29652 7140 31948
rect 7420 31332 7476 33182
rect 7644 33124 7700 34750
rect 7868 34354 7924 34860
rect 8092 34822 8148 34860
rect 7868 34302 7870 34354
rect 7922 34302 7924 34354
rect 7868 34290 7924 34302
rect 8316 34244 8372 35868
rect 8988 35588 9044 36204
rect 8988 35522 9044 35532
rect 8540 35252 8596 35262
rect 8316 34188 8484 34244
rect 8204 34020 8260 34030
rect 8316 34020 8372 34030
rect 8260 34018 8372 34020
rect 8260 33966 8318 34018
rect 8370 33966 8372 34018
rect 8260 33964 8372 33966
rect 7644 33068 7812 33124
rect 7420 31266 7476 31276
rect 7644 32900 7700 32910
rect 7532 30882 7588 30894
rect 7532 30830 7534 30882
rect 7586 30830 7588 30882
rect 7532 30548 7588 30830
rect 7532 30482 7588 30492
rect 7532 30100 7588 30110
rect 7644 30100 7700 32844
rect 7756 32788 7812 33068
rect 7756 32722 7812 32732
rect 8092 31668 8148 31678
rect 7980 31612 8092 31668
rect 7868 30212 7924 30222
rect 7868 30118 7924 30156
rect 7532 30098 7700 30100
rect 7532 30046 7534 30098
rect 7586 30046 7700 30098
rect 7532 30044 7700 30046
rect 7532 30034 7588 30044
rect 7532 29876 7588 29886
rect 7084 29650 7476 29652
rect 7084 29598 7086 29650
rect 7138 29598 7476 29650
rect 7084 29596 7476 29598
rect 7084 29586 7140 29596
rect 7420 29316 7476 29596
rect 7532 29538 7588 29820
rect 7532 29486 7534 29538
rect 7586 29486 7588 29538
rect 7532 29474 7588 29486
rect 7980 29426 8036 31612
rect 8092 31602 8148 31612
rect 7980 29374 7982 29426
rect 8034 29374 8036 29426
rect 7644 29316 7700 29326
rect 7420 29314 7700 29316
rect 7420 29262 7646 29314
rect 7698 29262 7700 29314
rect 7420 29260 7700 29262
rect 7644 29250 7700 29260
rect 7532 28756 7588 28766
rect 6972 28532 7028 28542
rect 6972 28530 7140 28532
rect 6972 28478 6974 28530
rect 7026 28478 7140 28530
rect 6972 28476 7140 28478
rect 6972 28466 7028 28476
rect 7084 28082 7140 28476
rect 7084 28030 7086 28082
rect 7138 28030 7140 28082
rect 7084 28018 7140 28030
rect 6972 27860 7028 27870
rect 6972 27766 7028 27804
rect 7308 26292 7364 26302
rect 6860 26290 7364 26292
rect 6860 26238 7310 26290
rect 7362 26238 7364 26290
rect 6860 26236 7364 26238
rect 7308 26226 7364 26236
rect 7084 26066 7140 26078
rect 7084 26014 7086 26066
rect 7138 26014 7140 26066
rect 7084 25620 7140 26014
rect 7308 25620 7364 25630
rect 7084 25564 7308 25620
rect 7308 25526 7364 25564
rect 7532 25508 7588 28700
rect 7980 28532 8036 29374
rect 7980 28466 8036 28476
rect 8092 29652 8148 29662
rect 7980 28084 8036 28094
rect 8092 28084 8148 29596
rect 7980 28082 8148 28084
rect 7980 28030 7982 28082
rect 8034 28030 8148 28082
rect 7980 28028 8148 28030
rect 7980 28018 8036 28028
rect 7756 27972 7812 27982
rect 7756 27858 7812 27916
rect 7756 27806 7758 27858
rect 7810 27806 7812 27858
rect 7756 27794 7812 27806
rect 8092 27860 8148 28028
rect 8092 27794 8148 27804
rect 8092 26964 8148 27002
rect 7868 26852 8148 26908
rect 8204 26908 8260 33964
rect 8316 33954 8372 33964
rect 8428 33796 8484 34188
rect 8540 34130 8596 35196
rect 8540 34078 8542 34130
rect 8594 34078 8596 34130
rect 8540 34066 8596 34078
rect 8652 34914 8708 34926
rect 8652 34862 8654 34914
rect 8706 34862 8708 34914
rect 8316 33740 8484 33796
rect 8316 33458 8372 33740
rect 8316 33406 8318 33458
rect 8370 33406 8372 33458
rect 8316 33394 8372 33406
rect 8428 33234 8484 33246
rect 8428 33182 8430 33234
rect 8482 33182 8484 33234
rect 8428 31444 8484 33182
rect 8540 32450 8596 32462
rect 8540 32398 8542 32450
rect 8594 32398 8596 32450
rect 8540 31780 8596 32398
rect 8652 32116 8708 34862
rect 8876 33906 8932 33918
rect 8876 33854 8878 33906
rect 8930 33854 8932 33906
rect 8876 32900 8932 33854
rect 8876 32834 8932 32844
rect 9100 32676 9156 40350
rect 9548 38388 9604 40796
rect 9548 38322 9604 38332
rect 9548 38052 9604 38062
rect 9436 38050 9604 38052
rect 9436 37998 9550 38050
rect 9602 37998 9604 38050
rect 9436 37996 9604 37998
rect 9212 37826 9268 37838
rect 9212 37774 9214 37826
rect 9266 37774 9268 37826
rect 9212 37604 9268 37774
rect 9212 37538 9268 37548
rect 9212 33348 9268 33358
rect 9212 33254 9268 33292
rect 9100 32610 9156 32620
rect 8988 32562 9044 32574
rect 8988 32510 8990 32562
rect 9042 32510 9044 32562
rect 8988 32452 9044 32510
rect 9212 32564 9268 32574
rect 8988 32396 9156 32452
rect 8652 32050 8708 32060
rect 9100 31892 9156 32396
rect 9100 31826 9156 31836
rect 8988 31780 9044 31790
rect 8540 31778 9044 31780
rect 8540 31726 8990 31778
rect 9042 31726 9044 31778
rect 8540 31724 9044 31726
rect 8428 31378 8484 31388
rect 8988 30996 9044 31724
rect 9100 31556 9156 31566
rect 9100 31218 9156 31500
rect 9100 31166 9102 31218
rect 9154 31166 9156 31218
rect 9100 31154 9156 31166
rect 8652 30882 8708 30894
rect 8652 30830 8654 30882
rect 8706 30830 8708 30882
rect 8652 30770 8708 30830
rect 8652 30718 8654 30770
rect 8706 30718 8708 30770
rect 8652 30706 8708 30718
rect 8428 30212 8484 30222
rect 8428 28084 8484 30156
rect 8316 28028 8484 28084
rect 8540 30100 8596 30110
rect 8540 29764 8596 30044
rect 8540 28082 8596 29708
rect 8540 28030 8542 28082
rect 8594 28030 8596 28082
rect 8316 27636 8372 28028
rect 8428 27860 8484 27870
rect 8540 27860 8596 28030
rect 8652 29540 8708 29550
rect 8652 28082 8708 29484
rect 8876 29426 8932 29438
rect 8876 29374 8878 29426
rect 8930 29374 8932 29426
rect 8876 28868 8932 29374
rect 8876 28802 8932 28812
rect 8652 28030 8654 28082
rect 8706 28030 8708 28082
rect 8652 28018 8708 28030
rect 8764 28084 8820 28094
rect 8764 27990 8820 28028
rect 8988 27970 9044 30940
rect 9100 30770 9156 30782
rect 9100 30718 9102 30770
rect 9154 30718 9156 30770
rect 9100 30210 9156 30718
rect 9212 30322 9268 32508
rect 9324 31778 9380 31790
rect 9324 31726 9326 31778
rect 9378 31726 9380 31778
rect 9324 30548 9380 31726
rect 9436 31556 9492 37996
rect 9548 37986 9604 37996
rect 9548 37380 9604 37390
rect 9548 37154 9604 37324
rect 9548 37102 9550 37154
rect 9602 37102 9604 37154
rect 9548 35028 9604 37102
rect 9660 35924 9716 40910
rect 9772 40516 9828 40526
rect 9772 40422 9828 40460
rect 9884 38668 9940 41020
rect 9996 40516 10052 41244
rect 9996 40402 10052 40460
rect 9996 40350 9998 40402
rect 10050 40350 10052 40402
rect 9996 40338 10052 40350
rect 9884 38612 10052 38668
rect 9772 38164 9828 38174
rect 9772 37378 9828 38108
rect 9996 38050 10052 38612
rect 9996 37998 9998 38050
rect 10050 37998 10052 38050
rect 9996 37986 10052 37998
rect 10220 38052 10276 42252
rect 10444 41972 10500 45614
rect 10668 45220 10724 45230
rect 10668 44996 10724 45164
rect 10668 44930 10724 44940
rect 10780 44548 10836 46060
rect 11116 46004 11172 46014
rect 10892 45892 10948 45902
rect 10892 45788 10948 45836
rect 10892 45736 10894 45788
rect 10946 45736 10948 45788
rect 10892 45724 10948 45736
rect 10668 44492 10836 44548
rect 10892 45556 10948 45566
rect 10556 44210 10612 44222
rect 10556 44158 10558 44210
rect 10610 44158 10612 44210
rect 10556 42644 10612 44158
rect 10556 42578 10612 42588
rect 10444 41906 10500 41916
rect 10556 41970 10612 41982
rect 10556 41918 10558 41970
rect 10610 41918 10612 41970
rect 10556 41860 10612 41918
rect 10668 41972 10724 44492
rect 10892 44436 10948 45500
rect 10780 44380 10948 44436
rect 10780 43428 10836 44380
rect 11004 44324 11060 44334
rect 11004 44230 11060 44268
rect 11116 43876 11172 45948
rect 11228 45556 11284 48188
rect 11340 48178 11396 48188
rect 11564 48242 11844 48244
rect 11564 48190 11790 48242
rect 11842 48190 11844 48242
rect 11564 48188 11844 48190
rect 11340 48020 11396 48030
rect 11340 46786 11396 47964
rect 11452 47012 11508 47022
rect 11564 47012 11620 48188
rect 11788 48178 11844 48188
rect 11508 46956 11620 47012
rect 11452 46946 11508 46956
rect 11340 46734 11342 46786
rect 11394 46734 11396 46786
rect 11340 46722 11396 46734
rect 11452 46676 11508 46686
rect 11452 46582 11508 46620
rect 11900 46004 11956 48412
rect 12124 48356 12180 48366
rect 12124 48262 12180 48300
rect 11900 45938 11956 45948
rect 12124 45890 12180 45902
rect 12124 45838 12126 45890
rect 12178 45838 12180 45890
rect 11228 45490 11284 45500
rect 11676 45780 11732 45790
rect 12124 45780 12180 45838
rect 11732 45724 12180 45780
rect 11228 45332 11284 45342
rect 11228 45238 11284 45276
rect 11340 44996 11396 45006
rect 11340 44322 11396 44940
rect 11340 44270 11342 44322
rect 11394 44270 11396 44322
rect 11340 44258 11396 44270
rect 11452 44994 11508 45006
rect 11452 44942 11454 44994
rect 11506 44942 11508 44994
rect 11116 43820 11284 43876
rect 11116 43652 11172 43662
rect 11116 43558 11172 43596
rect 10780 42754 10836 43372
rect 10892 43538 10948 43550
rect 10892 43486 10894 43538
rect 10946 43486 10948 43538
rect 10892 42868 10948 43486
rect 10892 42802 10948 42812
rect 10780 42702 10782 42754
rect 10834 42702 10836 42754
rect 10780 42690 10836 42702
rect 10892 42530 10948 42542
rect 10892 42478 10894 42530
rect 10946 42478 10948 42530
rect 10668 41916 10836 41972
rect 10612 41804 10724 41860
rect 10556 41794 10612 41804
rect 10444 40068 10500 40078
rect 10332 40012 10444 40068
rect 10332 38164 10388 40012
rect 10444 40002 10500 40012
rect 10668 39618 10724 41804
rect 10668 39566 10670 39618
rect 10722 39566 10724 39618
rect 10668 39554 10724 39566
rect 10780 39620 10836 41916
rect 10892 40068 10948 42478
rect 11228 42084 11284 43820
rect 11452 43764 11508 44942
rect 11564 44324 11620 44334
rect 11676 44324 11732 45724
rect 11564 44322 11732 44324
rect 11564 44270 11566 44322
rect 11618 44270 11732 44322
rect 11564 44268 11732 44270
rect 12012 45444 12068 45454
rect 11564 44258 11620 44268
rect 11452 43698 11508 43708
rect 11788 44098 11844 44110
rect 11788 44046 11790 44098
rect 11842 44046 11844 44098
rect 11340 42642 11396 42654
rect 11340 42590 11342 42642
rect 11394 42590 11396 42642
rect 11340 42532 11396 42590
rect 11340 42466 11396 42476
rect 11676 42644 11732 42654
rect 10892 40002 10948 40012
rect 11116 42082 11284 42084
rect 11116 42030 11230 42082
rect 11282 42030 11284 42082
rect 11116 42028 11284 42030
rect 11116 39732 11172 42028
rect 11228 42018 11284 42028
rect 11340 40290 11396 40302
rect 11340 40238 11342 40290
rect 11394 40238 11396 40290
rect 10780 38836 10836 39564
rect 10780 38770 10836 38780
rect 10892 39730 11172 39732
rect 10892 39678 11118 39730
rect 11170 39678 11172 39730
rect 10892 39676 11172 39678
rect 10332 38108 10500 38164
rect 10220 37996 10388 38052
rect 9772 37326 9774 37378
rect 9826 37326 9828 37378
rect 9772 37314 9828 37326
rect 9884 37266 9940 37278
rect 9884 37214 9886 37266
rect 9938 37214 9940 37266
rect 9660 35868 9828 35924
rect 9660 35700 9716 35710
rect 9660 35606 9716 35644
rect 9660 35028 9716 35038
rect 9548 34972 9660 35028
rect 9660 34962 9716 34972
rect 9772 34804 9828 35868
rect 9548 34748 9828 34804
rect 9548 31892 9604 34748
rect 9660 34580 9716 34590
rect 9660 34130 9716 34524
rect 9660 34078 9662 34130
rect 9714 34078 9716 34130
rect 9660 34066 9716 34078
rect 9660 33348 9716 33358
rect 9660 33254 9716 33292
rect 9548 31826 9604 31836
rect 9660 32900 9716 32910
rect 9660 31778 9716 32844
rect 9884 32564 9940 37214
rect 10108 37268 10164 37278
rect 10108 37174 10164 37212
rect 9996 36708 10052 36718
rect 10052 36652 10164 36708
rect 9996 36642 10052 36652
rect 9996 35924 10052 35934
rect 9996 35830 10052 35868
rect 9996 35252 10052 35262
rect 9996 35026 10052 35196
rect 9996 34974 9998 35026
rect 10050 34974 10052 35026
rect 9996 34962 10052 34974
rect 10108 34356 10164 36652
rect 10220 36372 10276 36382
rect 10220 35922 10276 36316
rect 10220 35870 10222 35922
rect 10274 35870 10276 35922
rect 10220 35858 10276 35870
rect 10332 35922 10388 37996
rect 10444 37268 10500 38108
rect 10892 37938 10948 39676
rect 11116 39666 11172 39676
rect 11228 40068 11284 40078
rect 11116 38836 11172 38846
rect 11116 38164 11172 38780
rect 11116 38070 11172 38108
rect 10892 37886 10894 37938
rect 10946 37886 10948 37938
rect 10892 37874 10948 37886
rect 10668 37826 10724 37838
rect 10668 37774 10670 37826
rect 10722 37774 10724 37826
rect 10668 37716 10724 37774
rect 10668 37650 10724 37660
rect 11116 37826 11172 37838
rect 11116 37774 11118 37826
rect 11170 37774 11172 37826
rect 11116 37716 11172 37774
rect 10556 37492 10612 37502
rect 10556 37398 10612 37436
rect 11116 37380 11172 37660
rect 11116 37314 11172 37324
rect 10444 37212 10612 37268
rect 10444 36372 10500 36382
rect 10444 36278 10500 36316
rect 10332 35870 10334 35922
rect 10386 35870 10388 35922
rect 10332 35858 10388 35870
rect 10444 35924 10500 35934
rect 10444 34916 10500 35868
rect 10108 34290 10164 34300
rect 10220 34914 10500 34916
rect 10220 34862 10446 34914
rect 10498 34862 10500 34914
rect 10220 34860 10500 34862
rect 10108 34018 10164 34030
rect 10108 33966 10110 34018
rect 10162 33966 10164 34018
rect 10108 33460 10164 33966
rect 10108 33366 10164 33404
rect 10220 32676 10276 34860
rect 10444 34850 10500 34860
rect 10556 34580 10612 37212
rect 10892 36372 10948 36382
rect 10668 35924 10724 35934
rect 10668 35830 10724 35868
rect 10892 34914 10948 36316
rect 10892 34862 10894 34914
rect 10946 34862 10948 34914
rect 10892 34850 10948 34862
rect 11004 34802 11060 34814
rect 11004 34750 11006 34802
rect 11058 34750 11060 34802
rect 10612 34524 10836 34580
rect 10556 34514 10612 34524
rect 10220 32610 10276 32620
rect 10444 34356 10500 34366
rect 10444 33908 10500 34300
rect 10556 34244 10612 34282
rect 10556 34178 10612 34188
rect 10668 34130 10724 34142
rect 10668 34078 10670 34130
rect 10722 34078 10724 34130
rect 10556 33908 10612 33918
rect 10444 33906 10612 33908
rect 10444 33854 10558 33906
rect 10610 33854 10612 33906
rect 10444 33852 10612 33854
rect 9884 32498 9940 32508
rect 10332 32564 10388 32574
rect 10332 32470 10388 32508
rect 9660 31726 9662 31778
rect 9714 31726 9716 31778
rect 9660 31714 9716 31726
rect 9436 31490 9492 31500
rect 9884 31556 9940 31566
rect 9324 30492 9604 30548
rect 9212 30270 9214 30322
rect 9266 30270 9268 30322
rect 9212 30258 9268 30270
rect 9100 30158 9102 30210
rect 9154 30158 9156 30210
rect 9100 29204 9156 30158
rect 9548 30100 9604 30492
rect 9884 30210 9940 31500
rect 10108 30996 10164 31006
rect 10108 30902 10164 30940
rect 9884 30158 9886 30210
rect 9938 30158 9940 30210
rect 9660 30100 9716 30110
rect 9548 30044 9660 30100
rect 9660 30006 9716 30044
rect 9772 29540 9828 29550
rect 9772 29446 9828 29484
rect 9660 29428 9716 29438
rect 9660 29334 9716 29372
rect 9884 29316 9940 30158
rect 10220 29428 10276 29438
rect 10444 29428 10500 33852
rect 10556 33842 10612 33852
rect 10668 33460 10724 34078
rect 10668 33394 10724 33404
rect 10780 32788 10836 34524
rect 11004 34356 11060 34750
rect 10220 29426 10500 29428
rect 10220 29374 10222 29426
rect 10274 29374 10500 29426
rect 10220 29372 10500 29374
rect 10556 32732 10836 32788
rect 10892 34300 11060 34356
rect 11116 34802 11172 34814
rect 11116 34750 11118 34802
rect 11170 34750 11172 34802
rect 10220 29362 10276 29372
rect 9772 29260 9940 29316
rect 9772 29204 9828 29260
rect 10220 29204 10276 29214
rect 9100 29138 9156 29148
rect 9660 29148 9828 29204
rect 10108 29202 10276 29204
rect 10108 29150 10222 29202
rect 10274 29150 10276 29202
rect 10108 29148 10276 29150
rect 8988 27918 8990 27970
rect 9042 27918 9044 27970
rect 8988 27906 9044 27918
rect 8540 27804 8932 27860
rect 8428 27766 8484 27804
rect 8316 27580 8484 27636
rect 8204 26852 8372 26908
rect 7644 26404 7700 26414
rect 7644 26310 7700 26348
rect 7868 26402 7924 26852
rect 7868 26350 7870 26402
rect 7922 26350 7924 26402
rect 7868 26338 7924 26350
rect 8204 26290 8260 26302
rect 8204 26238 8206 26290
rect 8258 26238 8260 26290
rect 7756 26068 7812 26078
rect 7756 25974 7812 26012
rect 8204 25620 8260 26238
rect 7644 25618 8260 25620
rect 7644 25566 8206 25618
rect 8258 25566 8260 25618
rect 7644 25564 8260 25566
rect 7644 25508 7700 25564
rect 8204 25554 8260 25564
rect 7420 25506 7700 25508
rect 7420 25454 7646 25506
rect 7698 25454 7700 25506
rect 7420 25452 7700 25454
rect 6860 25396 6916 25406
rect 7420 25396 7476 25452
rect 7644 25442 7700 25452
rect 6860 25394 7476 25396
rect 6860 25342 6862 25394
rect 6914 25342 7476 25394
rect 6860 25340 7476 25342
rect 6860 25330 6916 25340
rect 8316 23268 8372 26852
rect 8428 25620 8484 27580
rect 8876 27186 8932 27804
rect 9100 27748 9156 27758
rect 9100 27300 9156 27692
rect 8876 27134 8878 27186
rect 8930 27134 8932 27186
rect 8876 27122 8932 27134
rect 8988 27244 9156 27300
rect 8764 26178 8820 26190
rect 8764 26126 8766 26178
rect 8818 26126 8820 26178
rect 8540 25620 8596 25630
rect 8428 25618 8596 25620
rect 8428 25566 8542 25618
rect 8594 25566 8596 25618
rect 8428 25564 8596 25566
rect 8540 25554 8596 25564
rect 8764 24836 8820 26126
rect 8988 25506 9044 27244
rect 9212 27188 9268 27198
rect 9212 27094 9268 27132
rect 9100 27076 9156 27086
rect 9100 26982 9156 27020
rect 9324 26852 9380 26862
rect 9324 26758 9380 26796
rect 9548 26852 9604 26862
rect 9660 26852 9716 29148
rect 10108 28642 10164 29148
rect 10220 29138 10276 29148
rect 10556 29092 10612 32732
rect 10780 32564 10836 32574
rect 10668 32452 10724 32462
rect 10780 32452 10836 32508
rect 10668 32450 10836 32452
rect 10668 32398 10670 32450
rect 10722 32398 10836 32450
rect 10668 32396 10836 32398
rect 10668 32386 10724 32396
rect 10668 30100 10724 30110
rect 10780 30100 10836 32396
rect 10892 32340 10948 34300
rect 11116 34244 11172 34750
rect 11004 34188 11172 34244
rect 11004 33906 11060 34188
rect 11004 33854 11006 33906
rect 11058 33854 11060 33906
rect 11004 33842 11060 33854
rect 11116 34020 11172 34030
rect 11116 33684 11172 33964
rect 11116 33618 11172 33628
rect 10892 32274 10948 32284
rect 11004 31778 11060 31790
rect 11004 31726 11006 31778
rect 11058 31726 11060 31778
rect 10892 31444 10948 31454
rect 10892 31218 10948 31388
rect 10892 31166 10894 31218
rect 10946 31166 10948 31218
rect 10892 31154 10948 31166
rect 11004 31108 11060 31726
rect 11004 30994 11060 31052
rect 11228 30996 11284 40012
rect 11340 36036 11396 40238
rect 11564 39396 11620 39406
rect 11564 39302 11620 39340
rect 11676 38668 11732 42588
rect 11788 42084 11844 44046
rect 11788 42018 11844 42028
rect 11900 43764 11956 43774
rect 11900 41186 11956 43708
rect 12012 41410 12068 45388
rect 12348 44436 12404 50372
rect 12460 49364 12516 52332
rect 12796 52276 12852 52668
rect 12796 52182 12852 52220
rect 14588 52276 14644 54462
rect 14924 54514 14980 54526
rect 14924 54462 14926 54514
rect 14978 54462 14980 54514
rect 14924 53508 14980 54462
rect 15708 54516 15764 54526
rect 15708 54422 15764 54460
rect 15932 54516 15988 54526
rect 16156 54516 16212 55356
rect 16380 55346 16436 55356
rect 16828 55300 16884 55310
rect 16828 55206 16884 55244
rect 15932 54514 16212 54516
rect 15932 54462 15934 54514
rect 15986 54462 16212 54514
rect 15932 54460 16212 54462
rect 16380 54516 16436 54526
rect 16828 54516 16884 54526
rect 16380 54514 16548 54516
rect 16380 54462 16382 54514
rect 16434 54462 16548 54514
rect 16380 54460 16548 54462
rect 15932 54450 15988 54460
rect 15932 53844 15988 53854
rect 15820 53788 15932 53844
rect 15372 53508 15428 53518
rect 14924 53506 15428 53508
rect 14924 53454 15374 53506
rect 15426 53454 15428 53506
rect 14924 53452 15428 53454
rect 14588 52162 14644 52220
rect 14588 52110 14590 52162
rect 14642 52110 14644 52162
rect 14588 52098 14644 52110
rect 14812 52724 14868 52734
rect 14812 52162 14868 52668
rect 15148 52612 15204 53452
rect 15372 53060 15428 53452
rect 15372 52994 15428 53004
rect 15372 52834 15428 52846
rect 15372 52782 15374 52834
rect 15426 52782 15428 52834
rect 15372 52724 15428 52782
rect 15372 52658 15428 52668
rect 14812 52110 14814 52162
rect 14866 52110 14868 52162
rect 14812 52098 14868 52110
rect 15036 52556 15204 52612
rect 14700 51938 14756 51950
rect 14700 51886 14702 51938
rect 14754 51886 14756 51938
rect 14700 51716 14756 51886
rect 13916 51660 14756 51716
rect 13916 51490 13972 51660
rect 15036 51604 15092 52556
rect 15148 52332 15652 52388
rect 15148 52162 15204 52332
rect 15596 52274 15652 52332
rect 15596 52222 15598 52274
rect 15650 52222 15652 52274
rect 15596 52210 15652 52222
rect 15148 52110 15150 52162
rect 15202 52110 15204 52162
rect 15148 52098 15204 52110
rect 15708 52162 15764 52174
rect 15708 52110 15710 52162
rect 15762 52110 15764 52162
rect 15484 51940 15540 51950
rect 15484 51846 15540 51884
rect 15036 51538 15092 51548
rect 13916 51438 13918 51490
rect 13970 51438 13972 51490
rect 13916 51426 13972 51438
rect 13132 51380 13188 51390
rect 15708 51380 15764 52110
rect 15820 52164 15876 53788
rect 15932 53778 15988 53788
rect 15932 53506 15988 53518
rect 15932 53454 15934 53506
rect 15986 53454 15988 53506
rect 15932 53172 15988 53454
rect 16044 53396 16100 54460
rect 16380 54450 16436 54460
rect 16492 53844 16548 54460
rect 16604 53844 16660 53854
rect 16492 53788 16604 53844
rect 16380 53730 16436 53742
rect 16380 53678 16382 53730
rect 16434 53678 16436 53730
rect 16044 53340 16212 53396
rect 15932 53106 15988 53116
rect 16044 52164 16100 52174
rect 15820 52162 16100 52164
rect 15820 52110 16046 52162
rect 16098 52110 16100 52162
rect 15820 52108 16100 52110
rect 16044 52098 16100 52108
rect 15708 51324 16100 51380
rect 13132 51286 13188 51324
rect 15820 50820 15876 50830
rect 15820 50428 15876 50764
rect 15932 50706 15988 51324
rect 16044 51266 16100 51324
rect 16044 51214 16046 51266
rect 16098 51214 16100 51266
rect 16044 51202 16100 51214
rect 15932 50654 15934 50706
rect 15986 50654 15988 50706
rect 15932 50642 15988 50654
rect 16156 50428 16212 53340
rect 16380 53172 16436 53678
rect 16604 53618 16660 53788
rect 16604 53566 16606 53618
rect 16658 53566 16660 53618
rect 16604 53554 16660 53566
rect 16380 53106 16436 53116
rect 16716 52500 16772 52510
rect 16492 52276 16548 52286
rect 16492 51602 16548 52220
rect 16492 51550 16494 51602
rect 16546 51550 16548 51602
rect 16492 51538 16548 51550
rect 16604 51380 16660 51390
rect 16492 50708 16548 50718
rect 16604 50708 16660 51324
rect 16492 50706 16660 50708
rect 16492 50654 16494 50706
rect 16546 50654 16660 50706
rect 16492 50652 16660 50654
rect 16492 50642 16548 50652
rect 16716 50428 16772 52444
rect 16828 51940 16884 54460
rect 17276 54514 17332 54526
rect 17276 54462 17278 54514
rect 17330 54462 17332 54514
rect 17276 52276 17332 54462
rect 17276 52210 17332 52220
rect 16828 51874 16884 51884
rect 16828 51378 16884 51390
rect 16828 51326 16830 51378
rect 16882 51326 16884 51378
rect 16828 50820 16884 51326
rect 16828 50754 16884 50764
rect 17388 50820 17444 50830
rect 17388 50594 17444 50764
rect 17388 50542 17390 50594
rect 17442 50542 17444 50594
rect 17388 50530 17444 50542
rect 12572 50370 12628 50382
rect 15820 50372 15988 50428
rect 12572 50318 12574 50370
rect 12626 50318 12628 50370
rect 12572 49812 12628 50318
rect 14364 50036 14420 50046
rect 13132 49922 13188 49934
rect 13132 49870 13134 49922
rect 13186 49870 13188 49922
rect 12572 49746 12628 49756
rect 12908 49810 12964 49822
rect 12908 49758 12910 49810
rect 12962 49758 12964 49810
rect 12460 49138 12516 49308
rect 12908 49364 12964 49758
rect 13132 49812 13188 49870
rect 12908 49298 12964 49308
rect 13020 49476 13076 49486
rect 12460 49086 12462 49138
rect 12514 49086 12516 49138
rect 12460 49074 12516 49086
rect 12684 47908 12740 47918
rect 12740 47852 12852 47908
rect 12684 47842 12740 47852
rect 12796 47346 12852 47852
rect 12796 47294 12798 47346
rect 12850 47294 12852 47346
rect 12796 47282 12852 47294
rect 12572 44436 12628 44446
rect 12348 44434 12628 44436
rect 12348 44382 12574 44434
rect 12626 44382 12628 44434
rect 12348 44380 12628 44382
rect 12572 44370 12628 44380
rect 12796 44322 12852 44334
rect 12796 44270 12798 44322
rect 12850 44270 12852 44322
rect 12460 44210 12516 44222
rect 12460 44158 12462 44210
rect 12514 44158 12516 44210
rect 12236 43764 12292 43774
rect 12012 41358 12014 41410
rect 12066 41358 12068 41410
rect 12012 41346 12068 41358
rect 12124 43652 12180 43662
rect 12124 42082 12180 43596
rect 12236 43538 12292 43708
rect 12460 43652 12516 44158
rect 12796 44100 12852 44270
rect 12796 44034 12852 44044
rect 13020 43988 13076 49420
rect 13132 47908 13188 49756
rect 14364 49138 14420 49980
rect 15260 50036 15316 50046
rect 15260 49942 15316 49980
rect 14364 49086 14366 49138
rect 14418 49086 14420 49138
rect 13916 49028 13972 49038
rect 14140 49028 14196 49038
rect 13916 49026 14084 49028
rect 13916 48974 13918 49026
rect 13970 48974 14084 49026
rect 13916 48972 14084 48974
rect 13916 48962 13972 48972
rect 13468 48804 13524 48814
rect 13468 48802 13748 48804
rect 13468 48750 13470 48802
rect 13522 48750 13748 48802
rect 13468 48748 13748 48750
rect 13468 48738 13524 48748
rect 13580 48580 13636 48590
rect 13580 48242 13636 48524
rect 13580 48190 13582 48242
rect 13634 48190 13636 48242
rect 13580 48178 13636 48190
rect 13132 47842 13188 47852
rect 13356 48132 13412 48142
rect 12460 43586 12516 43596
rect 12908 43932 13076 43988
rect 13132 46788 13188 46798
rect 13356 46788 13412 48076
rect 13692 46900 13748 48748
rect 14028 48580 14084 48972
rect 14140 49026 14308 49028
rect 14140 48974 14142 49026
rect 14194 48974 14308 49026
rect 14140 48972 14308 48974
rect 14140 48962 14196 48972
rect 14028 48514 14084 48524
rect 14252 48580 14308 48972
rect 14364 48804 14420 49086
rect 14924 49698 14980 49710
rect 14924 49646 14926 49698
rect 14978 49646 14980 49698
rect 14364 48738 14420 48748
rect 14812 48804 14868 48814
rect 14924 48804 14980 49646
rect 15708 49700 15764 49710
rect 14812 48802 14980 48804
rect 14812 48750 14814 48802
rect 14866 48750 14980 48802
rect 14812 48748 14980 48750
rect 15036 49252 15092 49262
rect 14812 48580 14868 48748
rect 14252 48524 14868 48580
rect 14252 48356 14308 48524
rect 13804 48300 14308 48356
rect 14364 48356 14420 48366
rect 13804 48242 13860 48300
rect 13804 48190 13806 48242
rect 13858 48190 13860 48242
rect 13804 48178 13860 48190
rect 14028 48018 14084 48030
rect 14028 47966 14030 48018
rect 14082 47966 14084 48018
rect 14028 47346 14084 47966
rect 14028 47294 14030 47346
rect 14082 47294 14084 47346
rect 13692 46898 13972 46900
rect 13692 46846 13694 46898
rect 13746 46846 13972 46898
rect 13692 46844 13972 46846
rect 13692 46834 13748 46844
rect 12236 43486 12238 43538
rect 12290 43486 12292 43538
rect 12236 43474 12292 43486
rect 12348 43428 12404 43438
rect 12572 43428 12628 43438
rect 12348 43426 12516 43428
rect 12348 43374 12350 43426
rect 12402 43374 12516 43426
rect 12348 43372 12516 43374
rect 12348 43362 12404 43372
rect 12124 42030 12126 42082
rect 12178 42030 12180 42082
rect 11900 41134 11902 41186
rect 11954 41134 11956 41186
rect 11900 41122 11956 41134
rect 12124 41074 12180 42030
rect 12348 42644 12404 42654
rect 12124 41022 12126 41074
rect 12178 41022 12180 41074
rect 12124 41010 12180 41022
rect 12236 41970 12292 41982
rect 12236 41918 12238 41970
rect 12290 41918 12292 41970
rect 12236 40852 12292 41918
rect 11900 40796 12292 40852
rect 11788 40516 11844 40526
rect 11788 40422 11844 40460
rect 11788 39620 11844 39630
rect 11900 39620 11956 40796
rect 12348 40626 12404 42588
rect 12348 40574 12350 40626
rect 12402 40574 12404 40626
rect 12348 40562 12404 40574
rect 12012 40292 12068 40302
rect 12460 40292 12516 43372
rect 12572 43334 12628 43372
rect 12908 40740 12964 43932
rect 13020 43540 13076 43550
rect 13132 43540 13188 46732
rect 13020 43538 13188 43540
rect 13020 43486 13022 43538
rect 13074 43486 13188 43538
rect 13020 43484 13188 43486
rect 13244 46786 13412 46788
rect 13244 46734 13358 46786
rect 13410 46734 13412 46786
rect 13244 46732 13412 46734
rect 13020 43474 13076 43484
rect 12068 40236 12516 40292
rect 12572 40684 12964 40740
rect 13132 41524 13188 41534
rect 12012 40198 12068 40236
rect 11844 39564 11956 39620
rect 11788 39554 11844 39564
rect 11340 35970 11396 35980
rect 11452 38612 11732 38668
rect 11788 39060 11844 39070
rect 11788 38668 11844 39004
rect 12348 38724 12404 38762
rect 11788 38612 11956 38668
rect 12348 38658 12404 38668
rect 12572 38668 12628 40684
rect 13132 40628 13188 41468
rect 12684 40626 13188 40628
rect 12684 40574 13134 40626
rect 13186 40574 13188 40626
rect 12684 40572 13188 40574
rect 12684 39730 12740 40572
rect 13132 40562 13188 40572
rect 12684 39678 12686 39730
rect 12738 39678 12740 39730
rect 12684 39666 12740 39678
rect 12908 40402 12964 40414
rect 13244 40404 13300 46732
rect 13356 46722 13412 46732
rect 13916 45890 13972 46844
rect 14028 46788 14084 47294
rect 14028 46722 14084 46732
rect 14364 46562 14420 48300
rect 14476 48244 14532 48254
rect 14476 48150 14532 48188
rect 14812 47460 14868 48524
rect 14924 47460 14980 47470
rect 14812 47458 14980 47460
rect 14812 47406 14926 47458
rect 14978 47406 14980 47458
rect 14812 47404 14980 47406
rect 14812 46900 14868 47404
rect 14924 47394 14980 47404
rect 15036 47234 15092 49196
rect 15148 49026 15204 49038
rect 15148 48974 15150 49026
rect 15202 48974 15204 49026
rect 15148 48244 15204 48974
rect 15148 48178 15204 48188
rect 15372 49026 15428 49038
rect 15372 48974 15374 49026
rect 15426 48974 15428 49026
rect 15372 48916 15428 48974
rect 15372 48242 15428 48860
rect 15708 48354 15764 49644
rect 15932 49138 15988 50372
rect 16044 50372 16100 50382
rect 16156 50372 16436 50428
rect 16044 50278 16100 50316
rect 15932 49086 15934 49138
rect 15986 49086 15988 49138
rect 15932 49074 15988 49086
rect 16268 50036 16324 50046
rect 15708 48302 15710 48354
rect 15762 48302 15764 48354
rect 15708 48290 15764 48302
rect 15820 48804 15876 48814
rect 15372 48190 15374 48242
rect 15426 48190 15428 48242
rect 15372 48178 15428 48190
rect 15260 48132 15316 48142
rect 15260 48038 15316 48076
rect 15036 47182 15038 47234
rect 15090 47182 15092 47234
rect 15036 47170 15092 47182
rect 15260 47458 15316 47470
rect 15260 47406 15262 47458
rect 15314 47406 15316 47458
rect 15260 47012 15316 47406
rect 15372 47012 15428 47022
rect 14812 46834 14868 46844
rect 14924 46956 15372 47012
rect 14700 46676 14756 46686
rect 14924 46676 14980 46956
rect 15372 46946 15428 46956
rect 14700 46674 14980 46676
rect 14700 46622 14702 46674
rect 14754 46622 14980 46674
rect 14700 46620 14980 46622
rect 15036 46788 15092 46798
rect 15036 46674 15092 46732
rect 15708 46788 15764 46798
rect 15708 46694 15764 46732
rect 15036 46622 15038 46674
rect 15090 46622 15092 46674
rect 14700 46610 14756 46620
rect 15036 46610 15092 46622
rect 14364 46510 14366 46562
rect 14418 46510 14420 46562
rect 14364 46498 14420 46510
rect 15036 46452 15092 46462
rect 15036 46358 15092 46396
rect 14476 46228 14532 46238
rect 14476 46002 14532 46172
rect 14476 45950 14478 46002
rect 14530 45950 14532 46002
rect 14476 45938 14532 45950
rect 13916 45838 13918 45890
rect 13970 45838 13972 45890
rect 13916 45826 13972 45838
rect 14812 45220 14868 45230
rect 13692 45108 13748 45118
rect 13692 45014 13748 45052
rect 14364 45108 14420 45118
rect 14252 44996 14308 45006
rect 14140 44994 14308 44996
rect 14140 44942 14254 44994
rect 14306 44942 14308 44994
rect 14140 44940 14308 44942
rect 13692 44100 13748 44110
rect 13692 44006 13748 44044
rect 14028 43988 14084 43998
rect 13468 43540 13524 43550
rect 13468 42754 13524 43484
rect 13916 43540 13972 43550
rect 13916 43446 13972 43484
rect 13916 42868 13972 42878
rect 13468 42702 13470 42754
rect 13522 42702 13524 42754
rect 13468 42690 13524 42702
rect 13580 42866 13972 42868
rect 13580 42814 13918 42866
rect 13970 42814 13972 42866
rect 13580 42812 13972 42814
rect 13356 41858 13412 41870
rect 13356 41806 13358 41858
rect 13410 41806 13412 41858
rect 13356 41524 13412 41806
rect 13356 41458 13412 41468
rect 13580 40964 13636 42812
rect 13916 42802 13972 42812
rect 14028 42308 14084 43932
rect 14028 42242 14084 42252
rect 13916 42084 13972 42094
rect 13916 41412 13972 42028
rect 14140 41636 14196 44940
rect 14252 44930 14308 44940
rect 14364 44322 14420 45052
rect 14812 44434 14868 45164
rect 14812 44382 14814 44434
rect 14866 44382 14868 44434
rect 14812 44370 14868 44382
rect 15260 44772 15316 44782
rect 14364 44270 14366 44322
rect 14418 44270 14420 44322
rect 14364 44258 14420 44270
rect 15260 44322 15316 44716
rect 15260 44270 15262 44322
rect 15314 44270 15316 44322
rect 14476 43876 14532 43886
rect 14476 43426 14532 43820
rect 14476 43374 14478 43426
rect 14530 43374 14532 43426
rect 14364 42196 14420 42206
rect 14140 41580 14308 41636
rect 13804 41410 13972 41412
rect 13804 41358 13918 41410
rect 13970 41358 13972 41410
rect 13804 41356 13972 41358
rect 13692 41076 13748 41086
rect 13692 40982 13748 41020
rect 12908 40350 12910 40402
rect 12962 40350 12964 40402
rect 12908 39508 12964 40350
rect 13132 40348 13300 40404
rect 13468 40908 13636 40964
rect 13020 40292 13076 40302
rect 13020 40198 13076 40236
rect 12908 39442 12964 39452
rect 13020 39060 13076 39070
rect 13020 38966 13076 39004
rect 12796 38834 12852 38846
rect 12796 38782 12798 38834
rect 12850 38782 12852 38834
rect 12572 38612 12740 38668
rect 11452 38050 11508 38612
rect 11452 37998 11454 38050
rect 11506 37998 11508 38050
rect 11340 35140 11396 35150
rect 11340 34356 11396 35084
rect 11452 34804 11508 37998
rect 11788 38050 11844 38062
rect 11788 37998 11790 38050
rect 11842 37998 11844 38050
rect 11788 37492 11844 37998
rect 11900 38050 11956 38612
rect 12236 38276 12292 38286
rect 12236 38162 12292 38220
rect 12236 38110 12238 38162
rect 12290 38110 12292 38162
rect 12236 38098 12292 38110
rect 11900 37998 11902 38050
rect 11954 37998 11956 38050
rect 11900 37986 11956 37998
rect 12348 38052 12404 38062
rect 12684 38052 12740 38612
rect 12796 38276 12852 38782
rect 12796 38210 12852 38220
rect 12796 38052 12852 38062
rect 12348 38050 12852 38052
rect 12348 37998 12350 38050
rect 12402 37998 12798 38050
rect 12850 37998 12852 38050
rect 12348 37996 12852 37998
rect 12348 37986 12404 37996
rect 12124 37828 12180 37838
rect 12124 37734 12180 37772
rect 12348 37828 12404 37838
rect 11900 37492 11956 37502
rect 11788 37436 11900 37492
rect 11900 37266 11956 37436
rect 11900 37214 11902 37266
rect 11954 37214 11956 37266
rect 11900 37202 11956 37214
rect 12124 37380 12180 37390
rect 11788 37044 11844 37054
rect 11788 35922 11844 36988
rect 12124 36260 12180 37324
rect 12124 36194 12180 36204
rect 11788 35870 11790 35922
rect 11842 35870 11844 35922
rect 11564 35588 11620 35598
rect 11564 35586 11732 35588
rect 11564 35534 11566 35586
rect 11618 35534 11732 35586
rect 11564 35532 11732 35534
rect 11564 35522 11620 35532
rect 11564 35364 11620 35374
rect 11564 35138 11620 35308
rect 11564 35086 11566 35138
rect 11618 35086 11620 35138
rect 11564 35074 11620 35086
rect 11452 34738 11508 34748
rect 11676 34692 11732 35532
rect 11788 34916 11844 35870
rect 12012 35924 12068 35934
rect 12012 35830 12068 35868
rect 12124 35700 12180 35710
rect 12124 35606 12180 35644
rect 11788 34850 11844 34860
rect 12236 35140 12292 35150
rect 12236 34914 12292 35084
rect 12348 35138 12404 37772
rect 12348 35086 12350 35138
rect 12402 35086 12404 35138
rect 12348 35074 12404 35086
rect 12236 34862 12238 34914
rect 12290 34862 12292 34914
rect 12012 34692 12068 34702
rect 11676 34690 12068 34692
rect 11676 34638 12014 34690
rect 12066 34638 12068 34690
rect 11676 34636 12068 34638
rect 12012 34468 12068 34636
rect 12012 34402 12068 34412
rect 11564 34356 11620 34366
rect 11340 34354 11620 34356
rect 11340 34302 11566 34354
rect 11618 34302 11620 34354
rect 11340 34300 11620 34302
rect 11564 34290 11620 34300
rect 12236 34356 12292 34862
rect 12460 34356 12516 37996
rect 12796 37986 12852 37996
rect 13020 37716 13076 37726
rect 12572 37492 12628 37502
rect 13020 37492 13076 37660
rect 12628 37490 13076 37492
rect 12628 37438 13022 37490
rect 13074 37438 13076 37490
rect 12628 37436 13076 37438
rect 12572 37398 12628 37436
rect 13020 37426 13076 37436
rect 12908 36596 12964 36606
rect 13132 36596 13188 40348
rect 13356 38948 13412 38958
rect 13244 38892 13356 38948
rect 13244 38500 13300 38892
rect 13356 38882 13412 38892
rect 13468 38668 13524 40908
rect 13580 40740 13636 40750
rect 13580 40402 13636 40684
rect 13580 40350 13582 40402
rect 13634 40350 13636 40402
rect 13580 40338 13636 40350
rect 13468 38612 13748 38668
rect 13244 38444 13636 38500
rect 13580 38274 13636 38444
rect 13580 38222 13582 38274
rect 13634 38222 13636 38274
rect 13580 38210 13636 38222
rect 13692 38052 13748 38612
rect 13580 37996 13748 38052
rect 13468 37938 13524 37950
rect 13468 37886 13470 37938
rect 13522 37886 13524 37938
rect 13468 37044 13524 37886
rect 13468 36978 13524 36988
rect 13580 36820 13636 37996
rect 13692 37828 13748 37838
rect 13692 37734 13748 37772
rect 12572 36594 13188 36596
rect 12572 36542 12910 36594
rect 12962 36542 13188 36594
rect 12572 36540 13188 36542
rect 12572 36372 12628 36540
rect 12908 36530 12964 36540
rect 13132 36484 13188 36540
rect 13132 36418 13188 36428
rect 13468 36764 13636 36820
rect 12572 35922 12628 36316
rect 12572 35870 12574 35922
rect 12626 35870 12628 35922
rect 12572 35858 12628 35870
rect 13020 35700 13076 35710
rect 13020 35586 13076 35644
rect 13020 35534 13022 35586
rect 13074 35534 13076 35586
rect 12572 34916 12628 34926
rect 12572 34822 12628 34860
rect 12908 34692 12964 34702
rect 13020 34692 13076 35534
rect 12908 34690 13076 34692
rect 12908 34638 12910 34690
rect 12962 34638 13076 34690
rect 12908 34636 13076 34638
rect 13132 35140 13188 35150
rect 12908 34356 12964 34636
rect 12236 34290 12292 34300
rect 12348 34300 12516 34356
rect 12572 34300 12964 34356
rect 12012 34020 12068 34030
rect 12012 33926 12068 33964
rect 11676 33906 11732 33918
rect 11676 33854 11678 33906
rect 11730 33854 11732 33906
rect 11452 31668 11508 31678
rect 11452 31574 11508 31612
rect 11004 30942 11006 30994
rect 11058 30942 11060 30994
rect 11004 30930 11060 30942
rect 11116 30940 11284 30996
rect 11452 30996 11508 31006
rect 11508 30940 11620 30996
rect 10780 30044 10948 30100
rect 10668 29988 10724 30044
rect 10668 29986 10836 29988
rect 10668 29934 10670 29986
rect 10722 29934 10836 29986
rect 10668 29932 10836 29934
rect 10668 29922 10724 29932
rect 10108 28590 10110 28642
rect 10162 28590 10164 28642
rect 10108 28578 10164 28590
rect 10444 29036 10612 29092
rect 10668 29428 10724 29438
rect 10220 28532 10276 28542
rect 10220 28438 10276 28476
rect 10444 27972 10500 29036
rect 10556 28868 10612 28878
rect 10556 28642 10612 28812
rect 10668 28754 10724 29372
rect 10780 29092 10836 29932
rect 10780 29026 10836 29036
rect 10668 28702 10670 28754
rect 10722 28702 10724 28754
rect 10668 28690 10724 28702
rect 10556 28590 10558 28642
rect 10610 28590 10612 28642
rect 10556 28578 10612 28590
rect 10892 28532 10948 30044
rect 11004 29428 11060 29438
rect 11004 29334 11060 29372
rect 11004 28532 11060 28542
rect 10892 28530 11060 28532
rect 10892 28478 11006 28530
rect 11058 28478 11060 28530
rect 10892 28476 11060 28478
rect 10444 27860 10500 27916
rect 10780 28420 10836 28430
rect 10556 27860 10612 27870
rect 10444 27858 10612 27860
rect 10444 27806 10558 27858
rect 10610 27806 10612 27858
rect 10444 27804 10612 27806
rect 10556 27794 10612 27804
rect 9996 27748 10052 27758
rect 9996 27654 10052 27692
rect 10780 27412 10836 28364
rect 10780 27346 10836 27356
rect 10556 27188 10612 27198
rect 10892 27188 10948 28476
rect 11004 28420 11060 28476
rect 11004 28354 11060 28364
rect 10556 27186 10948 27188
rect 10556 27134 10558 27186
rect 10610 27134 10948 27186
rect 10556 27132 10948 27134
rect 9772 27074 9828 27086
rect 9772 27022 9774 27074
rect 9826 27022 9828 27074
rect 9772 26964 9828 27022
rect 10556 27076 10612 27132
rect 10556 27010 10612 27020
rect 10108 26964 10164 26974
rect 9772 26962 10164 26964
rect 9772 26910 10110 26962
rect 10162 26910 10164 26962
rect 9772 26908 10164 26910
rect 11116 26908 11172 30940
rect 11452 30930 11508 30940
rect 11564 30212 11620 30940
rect 11676 30324 11732 33854
rect 12124 33236 12180 33246
rect 12124 32562 12180 33180
rect 12348 33012 12404 34300
rect 12460 34132 12516 34142
rect 12572 34132 12628 34300
rect 13132 34244 13188 35084
rect 13468 35140 13524 36764
rect 13804 36708 13860 41356
rect 13916 41346 13972 41356
rect 14140 41186 14196 41198
rect 14140 41134 14142 41186
rect 14194 41134 14196 41186
rect 13916 40964 13972 40974
rect 13916 39060 13972 40908
rect 14140 40516 14196 41134
rect 14140 40450 14196 40460
rect 13916 38052 13972 39004
rect 14140 39620 14196 39630
rect 14028 38834 14084 38846
rect 14028 38782 14030 38834
rect 14082 38782 14084 38834
rect 14028 38276 14084 38782
rect 14140 38500 14196 39564
rect 14140 38434 14196 38444
rect 14028 38220 14196 38276
rect 14028 38052 14084 38062
rect 13916 38050 14084 38052
rect 13916 37998 14030 38050
rect 14082 37998 14084 38050
rect 13916 37996 14084 37998
rect 14028 37986 14084 37996
rect 14140 37940 14196 38220
rect 14140 37874 14196 37884
rect 13916 37826 13972 37838
rect 13916 37774 13918 37826
rect 13970 37774 13972 37826
rect 13916 37492 13972 37774
rect 13916 37426 13972 37436
rect 14252 37268 14308 41580
rect 14364 41410 14420 42140
rect 14364 41358 14366 41410
rect 14418 41358 14420 41410
rect 14364 41346 14420 41358
rect 14364 40404 14420 40414
rect 14364 40310 14420 40348
rect 14476 40180 14532 43374
rect 14812 40964 14868 40974
rect 14812 40962 14980 40964
rect 14812 40910 14814 40962
rect 14866 40910 14980 40962
rect 14812 40908 14980 40910
rect 14812 40898 14868 40908
rect 14700 40516 14756 40526
rect 14700 40404 14756 40460
rect 14812 40404 14868 40414
rect 14700 40402 14868 40404
rect 14700 40350 14814 40402
rect 14866 40350 14868 40402
rect 14700 40348 14868 40350
rect 14812 40338 14868 40348
rect 14028 37212 14308 37268
rect 14364 40124 14532 40180
rect 13804 36652 13972 36708
rect 13804 36484 13860 36494
rect 13804 36370 13860 36428
rect 13804 36318 13806 36370
rect 13858 36318 13860 36370
rect 13804 36306 13860 36318
rect 13468 35074 13524 35084
rect 13580 36148 13636 36158
rect 12908 34132 12964 34142
rect 12516 34076 12628 34132
rect 12684 34130 12964 34132
rect 12684 34078 12910 34130
rect 12962 34078 12964 34130
rect 12684 34076 12964 34078
rect 12460 34038 12516 34076
rect 12684 34020 12740 34076
rect 12908 34066 12964 34076
rect 12348 32946 12404 32956
rect 12572 33122 12628 33134
rect 12572 33070 12574 33122
rect 12626 33070 12628 33122
rect 12124 32510 12126 32562
rect 12178 32510 12180 32562
rect 12124 32498 12180 32510
rect 12460 32452 12516 32462
rect 12460 32358 12516 32396
rect 12124 32004 12180 32014
rect 12012 31948 12124 32004
rect 11900 30994 11956 31006
rect 11900 30942 11902 30994
rect 11954 30942 11956 30994
rect 11788 30324 11844 30334
rect 11676 30322 11844 30324
rect 11676 30270 11790 30322
rect 11842 30270 11844 30322
rect 11676 30268 11844 30270
rect 11788 30258 11844 30268
rect 11900 30212 11956 30942
rect 11564 30156 11732 30212
rect 11228 30100 11284 30110
rect 11284 30044 11396 30100
rect 11228 30006 11284 30044
rect 11228 29204 11284 29214
rect 11228 28642 11284 29148
rect 11228 28590 11230 28642
rect 11282 28590 11284 28642
rect 11228 28578 11284 28590
rect 10108 26852 10276 26908
rect 11116 26852 11284 26908
rect 9660 26796 9828 26852
rect 9548 26290 9604 26796
rect 9772 26628 9828 26796
rect 9660 26516 9716 26526
rect 9660 26422 9716 26460
rect 9772 26514 9828 26572
rect 9772 26462 9774 26514
rect 9826 26462 9828 26514
rect 9772 26450 9828 26462
rect 10108 26516 10164 26526
rect 9548 26238 9550 26290
rect 9602 26238 9604 26290
rect 9548 25732 9604 26238
rect 9548 25666 9604 25676
rect 9660 26292 9716 26302
rect 9660 25620 9716 26236
rect 10108 26290 10164 26460
rect 10220 26404 10276 26852
rect 10556 26628 10612 26638
rect 10556 26514 10612 26572
rect 10556 26462 10558 26514
rect 10610 26462 10612 26514
rect 10332 26404 10388 26414
rect 10220 26348 10332 26404
rect 10332 26338 10388 26348
rect 10108 26238 10110 26290
rect 10162 26238 10164 26290
rect 10108 26226 10164 26238
rect 10556 26180 10612 26462
rect 10556 26114 10612 26124
rect 11004 26516 11060 26526
rect 8988 25454 8990 25506
rect 9042 25454 9044 25506
rect 8988 25442 9044 25454
rect 9436 25508 9492 25518
rect 9436 25414 9492 25452
rect 9660 25506 9716 25564
rect 9660 25454 9662 25506
rect 9714 25454 9716 25506
rect 9660 25442 9716 25454
rect 10220 26068 10276 26078
rect 10220 25506 10276 26012
rect 11004 26068 11060 26460
rect 11004 26002 11060 26012
rect 10220 25454 10222 25506
rect 10274 25454 10276 25506
rect 10220 25442 10276 25454
rect 10444 25506 10500 25518
rect 10444 25454 10446 25506
rect 10498 25454 10500 25506
rect 9548 25396 9604 25406
rect 9548 25302 9604 25340
rect 10444 25396 10500 25454
rect 11004 25508 11060 25518
rect 11004 25414 11060 25452
rect 10444 25330 10500 25340
rect 10780 25396 10836 25406
rect 10780 25302 10836 25340
rect 8764 24770 8820 24780
rect 9884 25282 9940 25294
rect 9884 25230 9886 25282
rect 9938 25230 9940 25282
rect 9884 24052 9940 25230
rect 11228 25284 11284 26852
rect 11340 26290 11396 30044
rect 11676 30098 11732 30156
rect 11900 30146 11956 30156
rect 11676 30046 11678 30098
rect 11730 30046 11732 30098
rect 11676 30034 11732 30046
rect 12012 30100 12068 31948
rect 12124 31938 12180 31948
rect 12348 31220 12404 31230
rect 12348 31108 12404 31164
rect 12236 31106 12404 31108
rect 12236 31054 12350 31106
rect 12402 31054 12404 31106
rect 12236 31052 12404 31054
rect 11564 29986 11620 29998
rect 11564 29934 11566 29986
rect 11618 29934 11620 29986
rect 11564 29876 11620 29934
rect 11900 29988 11956 29998
rect 12012 29988 12068 30044
rect 11900 29986 12068 29988
rect 11900 29934 11902 29986
rect 11954 29934 12068 29986
rect 11900 29932 12068 29934
rect 12124 30098 12180 30110
rect 12124 30046 12126 30098
rect 12178 30046 12180 30098
rect 11900 29922 11956 29932
rect 11676 29876 11732 29886
rect 11564 29820 11676 29876
rect 11676 29650 11732 29820
rect 11676 29598 11678 29650
rect 11730 29598 11732 29650
rect 11676 29586 11732 29598
rect 12012 29764 12068 29774
rect 11788 29428 11844 29438
rect 11788 28754 11844 29372
rect 12012 29314 12068 29708
rect 12124 29540 12180 30046
rect 12124 29474 12180 29484
rect 12236 30100 12292 31052
rect 12348 31042 12404 31052
rect 12572 30324 12628 33070
rect 12684 31444 12740 33964
rect 13020 33796 13076 33806
rect 12908 33236 12964 33246
rect 12796 33180 12908 33236
rect 12796 31778 12852 33180
rect 12908 33142 12964 33180
rect 12796 31726 12798 31778
rect 12850 31726 12852 31778
rect 12796 31714 12852 31726
rect 12908 32900 12964 32910
rect 12908 31554 12964 32844
rect 12908 31502 12910 31554
rect 12962 31502 12964 31554
rect 12908 31490 12964 31502
rect 12684 31388 12852 31444
rect 12012 29262 12014 29314
rect 12066 29262 12068 29314
rect 12012 29250 12068 29262
rect 11788 28702 11790 28754
rect 11842 28702 11844 28754
rect 11788 28690 11844 28702
rect 12124 29204 12180 29214
rect 12124 28754 12180 29148
rect 12124 28702 12126 28754
rect 12178 28702 12180 28754
rect 12124 28690 12180 28702
rect 11452 28420 11508 28430
rect 11452 28082 11508 28364
rect 11452 28030 11454 28082
rect 11506 28030 11508 28082
rect 11452 27972 11508 28030
rect 12236 28084 12292 30044
rect 12348 30268 12628 30324
rect 12348 29092 12404 30268
rect 12684 30212 12740 30222
rect 12572 30100 12628 30110
rect 12572 30006 12628 30044
rect 12684 30098 12740 30156
rect 12684 30046 12686 30098
rect 12738 30046 12740 30098
rect 12684 29650 12740 30046
rect 12684 29598 12686 29650
rect 12738 29598 12740 29650
rect 12684 29586 12740 29598
rect 12460 29428 12516 29438
rect 12796 29428 12852 31388
rect 13020 30436 13076 33740
rect 13132 33572 13188 34188
rect 13468 34916 13524 34926
rect 13132 33516 13412 33572
rect 13132 33348 13188 33358
rect 13132 32004 13188 33292
rect 13244 33012 13300 33022
rect 13244 32562 13300 32956
rect 13244 32510 13246 32562
rect 13298 32510 13300 32562
rect 13244 32452 13300 32510
rect 13244 32386 13300 32396
rect 13356 32116 13412 33516
rect 13468 33570 13524 34860
rect 13468 33518 13470 33570
rect 13522 33518 13524 33570
rect 13468 32786 13524 33518
rect 13468 32734 13470 32786
rect 13522 32734 13524 32786
rect 13468 32722 13524 32734
rect 13580 32116 13636 36092
rect 13916 35924 13972 36652
rect 14028 36484 14084 37212
rect 14140 36708 14196 36718
rect 14364 36708 14420 40124
rect 14924 39618 14980 40908
rect 15148 40962 15204 40974
rect 15148 40910 15150 40962
rect 15202 40910 15204 40962
rect 15148 40516 15204 40910
rect 15148 40450 15204 40460
rect 15260 40404 15316 44270
rect 15708 44324 15764 44334
rect 15708 44230 15764 44268
rect 15484 43428 15540 43438
rect 15260 40338 15316 40348
rect 15372 40402 15428 40414
rect 15372 40350 15374 40402
rect 15426 40350 15428 40402
rect 15372 40292 15428 40350
rect 14924 39566 14926 39618
rect 14978 39566 14980 39618
rect 14924 39554 14980 39566
rect 15260 40180 15316 40190
rect 14700 39396 14756 39406
rect 14476 39394 14756 39396
rect 14476 39342 14702 39394
rect 14754 39342 14756 39394
rect 14476 39340 14756 39342
rect 14476 39060 14532 39340
rect 14700 39330 14756 39340
rect 15260 39060 15316 40124
rect 15372 39732 15428 40236
rect 15372 39666 15428 39676
rect 14476 38834 14532 39004
rect 15148 39058 15316 39060
rect 15148 39006 15262 39058
rect 15314 39006 15316 39058
rect 15148 39004 15316 39006
rect 14476 38782 14478 38834
rect 14530 38782 14532 38834
rect 14476 38770 14532 38782
rect 14812 38834 14868 38846
rect 14812 38782 14814 38834
rect 14866 38782 14868 38834
rect 14812 38612 14868 38782
rect 15036 38836 15092 38846
rect 15036 38742 15092 38780
rect 14476 38500 14532 38510
rect 14532 38444 14644 38500
rect 14476 38434 14532 38444
rect 14476 37940 14532 37950
rect 14476 37846 14532 37884
rect 14140 36614 14196 36652
rect 14252 36652 14420 36708
rect 14028 36428 14196 36484
rect 13916 35698 13972 35868
rect 13916 35646 13918 35698
rect 13970 35646 13972 35698
rect 13916 35634 13972 35646
rect 14028 36258 14084 36270
rect 14028 36206 14030 36258
rect 14082 36206 14084 36258
rect 13916 35028 13972 35038
rect 13692 34804 13748 34814
rect 13692 34710 13748 34748
rect 13916 34354 13972 34972
rect 13916 34302 13918 34354
rect 13970 34302 13972 34354
rect 13916 34290 13972 34302
rect 14028 33796 14084 36206
rect 14028 33730 14084 33740
rect 14140 34130 14196 36428
rect 14140 34078 14142 34130
rect 14194 34078 14196 34130
rect 13916 33570 13972 33582
rect 13916 33518 13918 33570
rect 13970 33518 13972 33570
rect 13692 33122 13748 33134
rect 13692 33070 13694 33122
rect 13746 33070 13748 33122
rect 13692 33012 13748 33070
rect 13692 32946 13748 32956
rect 13132 31938 13188 31948
rect 13244 32060 13412 32116
rect 13468 32060 13636 32116
rect 13692 32452 13748 32462
rect 12908 30380 13076 30436
rect 13132 30884 13188 30894
rect 12908 30210 12964 30380
rect 12908 30158 12910 30210
rect 12962 30158 12964 30210
rect 12908 30146 12964 30158
rect 13020 30100 13076 30110
rect 12460 29426 12964 29428
rect 12460 29374 12462 29426
rect 12514 29374 12964 29426
rect 12460 29372 12964 29374
rect 12460 29362 12516 29372
rect 12684 29204 12740 29214
rect 12684 29202 12852 29204
rect 12684 29150 12686 29202
rect 12738 29150 12852 29202
rect 12684 29148 12852 29150
rect 12684 29138 12740 29148
rect 12404 29036 12516 29092
rect 12348 29026 12404 29036
rect 12236 28018 12292 28028
rect 11452 27906 11508 27916
rect 12012 27972 12068 27982
rect 12012 27636 12068 27916
rect 12348 27970 12404 27982
rect 12348 27918 12350 27970
rect 12402 27918 12404 27970
rect 12124 27860 12180 27870
rect 12124 27766 12180 27804
rect 12012 27580 12292 27636
rect 12124 26964 12180 27002
rect 12124 26898 12180 26908
rect 11340 26238 11342 26290
rect 11394 26238 11396 26290
rect 11340 26226 11396 26238
rect 11788 26852 11844 26862
rect 11788 25506 11844 26796
rect 11900 26292 11956 26302
rect 11900 26198 11956 26236
rect 12236 26290 12292 27580
rect 12236 26238 12238 26290
rect 12290 26238 12292 26290
rect 12236 26226 12292 26238
rect 12348 27076 12404 27918
rect 11788 25454 11790 25506
rect 11842 25454 11844 25506
rect 11788 25442 11844 25454
rect 11900 25508 11956 25518
rect 11900 25414 11956 25452
rect 12348 25506 12404 27020
rect 12348 25454 12350 25506
rect 12402 25454 12404 25506
rect 11228 24946 11284 25228
rect 11228 24894 11230 24946
rect 11282 24894 11284 24946
rect 11228 24882 11284 24894
rect 11340 25282 11396 25294
rect 11340 25230 11342 25282
rect 11394 25230 11396 25282
rect 9884 23986 9940 23996
rect 11340 23604 11396 25230
rect 12012 25284 12068 25294
rect 12012 25190 12068 25228
rect 11676 24948 11732 24958
rect 11676 24854 11732 24892
rect 12348 24948 12404 25454
rect 12348 24882 12404 24892
rect 12460 27188 12516 29036
rect 12684 28756 12740 28766
rect 12684 28662 12740 28700
rect 11676 24612 11732 24622
rect 11676 24050 11732 24556
rect 11676 23998 11678 24050
rect 11730 23998 11732 24050
rect 11676 23986 11732 23998
rect 12460 24050 12516 27132
rect 12572 28084 12628 28094
rect 12572 27186 12628 28028
rect 12572 27134 12574 27186
rect 12626 27134 12628 27186
rect 12572 27122 12628 27134
rect 12796 26740 12852 29148
rect 12908 26908 12964 29372
rect 13020 28082 13076 30044
rect 13132 29428 13188 30828
rect 13244 29428 13300 32060
rect 13468 31948 13524 32060
rect 13356 31892 13524 31948
rect 13580 31892 13636 31902
rect 13356 31332 13412 31892
rect 13356 31266 13412 31276
rect 13468 31778 13524 31790
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31220 13524 31726
rect 13468 31154 13524 31164
rect 13580 30210 13636 31836
rect 13692 31218 13748 32396
rect 13692 31166 13694 31218
rect 13746 31166 13748 31218
rect 13692 31154 13748 31166
rect 13804 32004 13860 32014
rect 13580 30158 13582 30210
rect 13634 30158 13636 30210
rect 13580 30146 13636 30158
rect 13804 29876 13860 31948
rect 13916 31668 13972 33518
rect 14140 33570 14196 34078
rect 14140 33518 14142 33570
rect 14194 33518 14196 33570
rect 14140 33506 14196 33518
rect 14028 33458 14084 33470
rect 14028 33406 14030 33458
rect 14082 33406 14084 33458
rect 14028 32900 14084 33406
rect 14140 33124 14196 33134
rect 14140 33030 14196 33068
rect 14028 32844 14196 32900
rect 14028 32676 14084 32714
rect 14028 32610 14084 32620
rect 14028 32452 14084 32462
rect 14028 31778 14084 32396
rect 14028 31726 14030 31778
rect 14082 31726 14084 31778
rect 14028 31714 14084 31726
rect 13916 31106 13972 31612
rect 14140 31556 14196 32844
rect 13916 31054 13918 31106
rect 13970 31054 13972 31106
rect 13916 31042 13972 31054
rect 14028 31500 14196 31556
rect 14028 30772 14084 31500
rect 14140 31332 14196 31342
rect 14140 31218 14196 31276
rect 14140 31166 14142 31218
rect 14194 31166 14196 31218
rect 14140 31154 14196 31166
rect 14252 31220 14308 36652
rect 14364 36484 14420 36494
rect 14364 36390 14420 36428
rect 14364 35586 14420 35598
rect 14364 35534 14366 35586
rect 14418 35534 14420 35586
rect 14364 34468 14420 35534
rect 14588 34468 14644 38444
rect 14812 36036 14868 38556
rect 15148 38162 15204 39004
rect 15260 38994 15316 39004
rect 15484 38946 15540 43372
rect 15708 41076 15764 41086
rect 15708 40982 15764 41020
rect 15820 40514 15876 48748
rect 16156 48804 16212 48814
rect 16156 48710 16212 48748
rect 16044 48692 16100 48702
rect 15932 48244 15988 48254
rect 15932 45890 15988 48188
rect 16044 46676 16100 48636
rect 16268 48468 16324 49980
rect 16380 48914 16436 50372
rect 16604 50372 16772 50428
rect 17500 50428 17556 56140
rect 19180 56194 19236 56206
rect 19180 56142 19182 56194
rect 19234 56142 19236 56194
rect 18508 55412 18564 55422
rect 17724 55300 17780 55310
rect 17724 55206 17780 55244
rect 18396 55188 18452 55198
rect 17836 55186 18452 55188
rect 17836 55134 18398 55186
rect 18450 55134 18452 55186
rect 17836 55132 18452 55134
rect 17836 54852 17892 55132
rect 18396 55122 18452 55132
rect 17612 54796 17892 54852
rect 17612 54738 17668 54796
rect 17612 54686 17614 54738
rect 17666 54686 17668 54738
rect 17612 54674 17668 54686
rect 18508 54738 18564 55356
rect 18508 54686 18510 54738
rect 18562 54686 18564 54738
rect 18508 54674 18564 54686
rect 18732 55300 18788 55310
rect 17612 54514 17668 54526
rect 17612 54462 17614 54514
rect 17666 54462 17668 54514
rect 17612 53732 17668 54462
rect 17836 54516 17892 54526
rect 17836 54422 17892 54460
rect 18284 54514 18340 54526
rect 18284 54462 18286 54514
rect 18338 54462 18340 54514
rect 18284 54404 18340 54462
rect 18396 54516 18452 54526
rect 18396 54422 18452 54460
rect 18284 54338 18340 54348
rect 17612 53508 17668 53676
rect 18172 53732 18228 53742
rect 18172 53638 18228 53676
rect 17612 53442 17668 53452
rect 17948 52946 18004 52958
rect 17948 52894 17950 52946
rect 18002 52894 18004 52946
rect 17836 52274 17892 52286
rect 17836 52222 17838 52274
rect 17890 52222 17892 52274
rect 17724 50596 17780 50606
rect 17724 50482 17780 50540
rect 17724 50430 17726 50482
rect 17778 50430 17780 50482
rect 17500 50372 17668 50428
rect 17724 50418 17780 50430
rect 17836 50428 17892 52222
rect 17948 52276 18004 52894
rect 18396 52946 18452 52958
rect 18396 52894 18398 52946
rect 18450 52894 18452 52946
rect 18172 52836 18228 52846
rect 18172 52742 18228 52780
rect 18396 52388 18452 52894
rect 18396 52322 18452 52332
rect 18508 52946 18564 52958
rect 18508 52894 18510 52946
rect 18562 52894 18564 52946
rect 17948 52210 18004 52220
rect 18508 52164 18564 52894
rect 18284 52108 18564 52164
rect 18172 51940 18228 51950
rect 18172 50596 18228 51884
rect 18284 50706 18340 52108
rect 18732 51490 18788 55244
rect 18732 51438 18734 51490
rect 18786 51438 18788 51490
rect 18732 51380 18788 51438
rect 18732 51314 18788 51324
rect 18844 54514 18900 54526
rect 18844 54462 18846 54514
rect 18898 54462 18900 54514
rect 18844 53844 18900 54462
rect 18284 50654 18286 50706
rect 18338 50654 18340 50706
rect 18284 50642 18340 50654
rect 18172 50530 18228 50540
rect 18844 50594 18900 53788
rect 19068 52834 19124 52846
rect 19068 52782 19070 52834
rect 19122 52782 19124 52834
rect 19068 52612 19124 52782
rect 19068 52388 19124 52556
rect 19068 52322 19124 52332
rect 18844 50542 18846 50594
rect 18898 50542 18900 50594
rect 18844 50530 18900 50542
rect 18396 50482 18452 50494
rect 18396 50430 18398 50482
rect 18450 50430 18452 50482
rect 18396 50428 18452 50430
rect 19180 50428 19236 56142
rect 20860 56196 20916 56252
rect 23100 56420 23156 59200
rect 25340 56420 25396 59200
rect 23100 56364 23604 56420
rect 23100 56306 23156 56364
rect 23100 56254 23102 56306
rect 23154 56254 23156 56306
rect 23100 56242 23156 56254
rect 21084 56196 21140 56206
rect 21420 56196 21476 56206
rect 20860 56194 21140 56196
rect 20860 56142 21086 56194
rect 21138 56142 21140 56194
rect 20860 56140 21140 56142
rect 21084 56130 21140 56140
rect 21308 56194 21476 56196
rect 21308 56142 21422 56194
rect 21474 56142 21476 56194
rect 21308 56140 21476 56142
rect 20524 55412 20580 55422
rect 20524 55318 20580 55356
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20972 54516 21028 54526
rect 20748 54514 21028 54516
rect 20748 54462 20974 54514
rect 21026 54462 21028 54514
rect 20748 54460 21028 54462
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19964 52836 20020 52846
rect 19964 52274 20020 52780
rect 19964 52222 19966 52274
rect 20018 52222 20020 52274
rect 19964 52210 20020 52222
rect 20748 52276 20804 54460
rect 20972 54450 21028 54460
rect 20748 52162 20804 52220
rect 20748 52110 20750 52162
rect 20802 52110 20804 52162
rect 20748 52098 20804 52110
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 17836 50372 18452 50428
rect 16604 50036 16660 50372
rect 16604 49970 16660 49980
rect 16492 49252 16548 49262
rect 17612 49252 17668 50372
rect 18396 49924 18452 50372
rect 18396 49858 18452 49868
rect 19068 50372 19236 50428
rect 21308 50428 21364 56140
rect 21420 56130 21476 56140
rect 23324 56194 23380 56206
rect 23324 56142 23326 56194
rect 23378 56142 23380 56194
rect 23324 55748 23380 56142
rect 23548 56082 23604 56364
rect 25340 56364 25844 56420
rect 25340 56306 25396 56364
rect 25340 56254 25342 56306
rect 25394 56254 25396 56306
rect 25340 56242 25396 56254
rect 23548 56030 23550 56082
rect 23602 56030 23604 56082
rect 23548 56018 23604 56030
rect 25564 56194 25620 56206
rect 25564 56142 25566 56194
rect 25618 56142 25620 56194
rect 22988 55692 23380 55748
rect 21420 55300 21476 55310
rect 21420 55206 21476 55244
rect 22988 55298 23044 55692
rect 22988 55246 22990 55298
rect 23042 55246 23044 55298
rect 22988 55234 23044 55246
rect 23324 55412 23380 55422
rect 22652 55076 22708 55086
rect 21756 54402 21812 54414
rect 21756 54350 21758 54402
rect 21810 54350 21812 54402
rect 21756 53732 21812 54350
rect 21756 53666 21812 53676
rect 21980 53844 22036 53854
rect 21980 53730 22036 53788
rect 22652 53844 22708 55020
rect 22876 55074 22932 55086
rect 22876 55022 22878 55074
rect 22930 55022 22932 55074
rect 22876 54516 22932 55022
rect 21980 53678 21982 53730
rect 22034 53678 22036 53730
rect 21980 53666 22036 53678
rect 22428 53732 22484 53742
rect 22428 53638 22484 53676
rect 22652 53730 22708 53788
rect 22652 53678 22654 53730
rect 22706 53678 22708 53730
rect 22652 53666 22708 53678
rect 22764 54460 22876 54516
rect 22316 53618 22372 53630
rect 22316 53566 22318 53618
rect 22370 53566 22372 53618
rect 22316 53508 22372 53566
rect 22316 52948 22372 53452
rect 22764 53060 22820 54460
rect 22876 54450 22932 54460
rect 22876 53844 22932 53854
rect 22876 53730 22932 53788
rect 22876 53678 22878 53730
rect 22930 53678 22932 53730
rect 22876 53666 22932 53678
rect 22764 52966 22820 53004
rect 21980 52946 22372 52948
rect 21980 52894 22318 52946
rect 22370 52894 22372 52946
rect 21980 52892 22372 52894
rect 21420 52276 21476 52286
rect 21420 50594 21476 52220
rect 21420 50542 21422 50594
rect 21474 50542 21476 50594
rect 21420 50530 21476 50542
rect 21980 50428 22036 52892
rect 22316 52882 22372 52892
rect 22988 52948 23044 52958
rect 22988 52946 23268 52948
rect 22988 52894 22990 52946
rect 23042 52894 23268 52946
rect 22988 52892 23268 52894
rect 22988 52882 23044 52892
rect 22540 52834 22596 52846
rect 22540 52782 22542 52834
rect 22594 52782 22596 52834
rect 22092 52276 22148 52286
rect 22092 52182 22148 52220
rect 22540 51604 22596 52782
rect 23100 52276 23156 52286
rect 23100 51604 23156 52220
rect 22092 51548 22596 51604
rect 22652 51602 23156 51604
rect 22652 51550 23102 51602
rect 23154 51550 23156 51602
rect 22652 51548 23156 51550
rect 22092 50706 22148 51548
rect 22652 51378 22708 51548
rect 23100 51538 23156 51548
rect 22652 51326 22654 51378
rect 22706 51326 22708 51378
rect 22652 51314 22708 51326
rect 22092 50654 22094 50706
rect 22146 50654 22148 50706
rect 22092 50642 22148 50654
rect 23212 50484 23268 52892
rect 21308 50372 21476 50428
rect 21980 50372 22820 50428
rect 23212 50418 23268 50428
rect 16492 49026 16548 49196
rect 16492 48974 16494 49026
rect 16546 48974 16548 49026
rect 16492 48962 16548 48974
rect 17276 49196 17668 49252
rect 16380 48862 16382 48914
rect 16434 48862 16436 48914
rect 16380 48850 16436 48862
rect 16716 48468 16772 48478
rect 16156 48466 16772 48468
rect 16156 48414 16270 48466
rect 16322 48414 16718 48466
rect 16770 48414 16772 48466
rect 16156 48412 16772 48414
rect 16156 47012 16212 48412
rect 16268 48402 16324 48412
rect 16716 48402 16772 48412
rect 17164 47460 17220 47470
rect 17164 47366 17220 47404
rect 17276 47346 17332 49196
rect 17612 49140 17668 49196
rect 17612 49084 18116 49140
rect 17500 49028 17556 49038
rect 17500 48354 17556 48972
rect 17612 48914 17668 49084
rect 18060 49026 18116 49084
rect 18060 48974 18062 49026
rect 18114 48974 18116 49026
rect 17612 48862 17614 48914
rect 17666 48862 17668 48914
rect 17612 48850 17668 48862
rect 17836 48916 17892 48926
rect 17836 48822 17892 48860
rect 17500 48302 17502 48354
rect 17554 48302 17556 48354
rect 17500 48290 17556 48302
rect 17948 48466 18004 48478
rect 17948 48414 17950 48466
rect 18002 48414 18004 48466
rect 17388 48018 17444 48030
rect 17388 47966 17390 48018
rect 17442 47966 17444 48018
rect 17388 47460 17444 47966
rect 17388 47394 17444 47404
rect 17276 47294 17278 47346
rect 17330 47294 17332 47346
rect 17276 47282 17332 47294
rect 16156 46898 16212 46956
rect 16156 46846 16158 46898
rect 16210 46846 16212 46898
rect 16156 46834 16212 46846
rect 16492 47234 16548 47246
rect 17500 47236 17556 47246
rect 16492 47182 16494 47234
rect 16546 47182 16548 47234
rect 16492 46788 16548 47182
rect 16492 46722 16548 46732
rect 17388 47234 17556 47236
rect 17388 47182 17502 47234
rect 17554 47182 17556 47234
rect 17388 47180 17556 47182
rect 16044 46620 16212 46676
rect 15932 45838 15934 45890
rect 15986 45838 15988 45890
rect 15932 45826 15988 45838
rect 16156 45778 16212 46620
rect 16380 46004 16436 46014
rect 16380 45890 16436 45948
rect 16380 45838 16382 45890
rect 16434 45838 16436 45890
rect 16380 45826 16436 45838
rect 16716 45892 16772 45902
rect 17276 45892 17332 45902
rect 16716 45890 17276 45892
rect 16716 45838 16718 45890
rect 16770 45838 17276 45890
rect 16716 45836 17276 45838
rect 16716 45826 16772 45836
rect 17276 45798 17332 45836
rect 16156 45726 16158 45778
rect 16210 45726 16212 45778
rect 16156 45714 16212 45726
rect 16044 45666 16100 45678
rect 16044 45614 16046 45666
rect 16098 45614 16100 45666
rect 16044 44436 16100 45614
rect 17276 45108 17332 45118
rect 17276 44546 17332 45052
rect 17276 44494 17278 44546
rect 17330 44494 17332 44546
rect 17276 44482 17332 44494
rect 16156 44436 16212 44446
rect 16044 44434 16212 44436
rect 16044 44382 16158 44434
rect 16210 44382 16212 44434
rect 16044 44380 16212 44382
rect 16156 44370 16212 44380
rect 16380 44322 16436 44334
rect 16380 44270 16382 44322
rect 16434 44270 16436 44322
rect 16380 43764 16436 44270
rect 16604 44322 16660 44334
rect 16604 44270 16606 44322
rect 16658 44270 16660 44322
rect 16604 43988 16660 44270
rect 16828 44324 16884 44334
rect 16828 44230 16884 44268
rect 16604 43922 16660 43932
rect 16380 43698 16436 43708
rect 17388 43650 17444 47180
rect 17500 47170 17556 47180
rect 17724 46004 17780 46014
rect 17724 45910 17780 45948
rect 17948 45780 18004 48414
rect 18060 48242 18116 48974
rect 18060 48190 18062 48242
rect 18114 48190 18116 48242
rect 18060 48178 18116 48190
rect 18284 49028 18340 49038
rect 18284 48130 18340 48972
rect 19068 49028 19124 50372
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20524 49252 20580 49262
rect 19068 48934 19124 48972
rect 19180 49138 19236 49150
rect 19180 49086 19182 49138
rect 19234 49086 19236 49138
rect 18396 48804 18452 48814
rect 18844 48804 18900 48814
rect 18396 48802 18900 48804
rect 18396 48750 18398 48802
rect 18450 48750 18846 48802
rect 18898 48750 18900 48802
rect 18396 48748 18900 48750
rect 18396 48738 18452 48748
rect 18284 48078 18286 48130
rect 18338 48078 18340 48130
rect 18284 48066 18340 48078
rect 18508 48580 18564 48590
rect 18284 47458 18340 47470
rect 18284 47406 18286 47458
rect 18338 47406 18340 47458
rect 17612 44436 17668 44446
rect 17612 44342 17668 44380
rect 17948 44212 18004 45724
rect 18172 47348 18228 47358
rect 18060 44212 18116 44222
rect 17948 44210 18116 44212
rect 17948 44158 18062 44210
rect 18114 44158 18116 44210
rect 17948 44156 18116 44158
rect 18060 44146 18116 44156
rect 17500 43764 17556 43774
rect 17500 43670 17556 43708
rect 18060 43764 18116 43774
rect 17388 43598 17390 43650
rect 17442 43598 17444 43650
rect 17388 43586 17444 43598
rect 17612 43652 17668 43662
rect 17612 43558 17668 43596
rect 17724 43650 17780 43662
rect 17724 43598 17726 43650
rect 17778 43598 17780 43650
rect 15820 40462 15822 40514
rect 15874 40462 15876 40514
rect 15820 40450 15876 40462
rect 15932 43540 15988 43550
rect 15484 38894 15486 38946
rect 15538 38894 15540 38946
rect 15372 38612 15428 38622
rect 15148 38110 15150 38162
rect 15202 38110 15204 38162
rect 15148 38098 15204 38110
rect 15260 38610 15428 38612
rect 15260 38558 15374 38610
rect 15426 38558 15428 38610
rect 15260 38556 15428 38558
rect 15036 38050 15092 38062
rect 15036 37998 15038 38050
rect 15090 37998 15092 38050
rect 15036 37716 15092 37998
rect 15036 37650 15092 37660
rect 15036 37268 15092 37278
rect 15260 37268 15316 38556
rect 15372 38546 15428 38556
rect 15372 37268 15428 37278
rect 15260 37266 15428 37268
rect 15260 37214 15374 37266
rect 15426 37214 15428 37266
rect 15260 37212 15428 37214
rect 14924 37154 14980 37166
rect 14924 37102 14926 37154
rect 14978 37102 14980 37154
rect 14924 36708 14980 37102
rect 14924 36642 14980 36652
rect 14812 35980 14980 36036
rect 14812 35812 14868 35822
rect 14812 35718 14868 35756
rect 14700 35698 14756 35710
rect 14700 35646 14702 35698
rect 14754 35646 14756 35698
rect 14700 35252 14756 35646
rect 14700 35186 14756 35196
rect 14812 35028 14868 35038
rect 14924 35028 14980 35980
rect 15036 35922 15092 37212
rect 15372 37202 15428 37212
rect 15148 37044 15204 37054
rect 15148 36950 15204 36988
rect 15484 36820 15540 38894
rect 15596 40404 15652 40414
rect 15596 38050 15652 40348
rect 15596 37998 15598 38050
rect 15650 37998 15652 38050
rect 15596 37986 15652 37998
rect 15708 39508 15764 39518
rect 15708 37156 15764 39452
rect 15820 37828 15876 37838
rect 15820 37734 15876 37772
rect 15820 37492 15876 37502
rect 15932 37492 15988 43484
rect 17724 43428 17780 43598
rect 17724 43362 17780 43372
rect 17836 43650 17892 43662
rect 17836 43598 17838 43650
rect 17890 43598 17892 43650
rect 17836 43204 17892 43598
rect 17500 43148 17892 43204
rect 16716 42196 16772 42206
rect 16716 42102 16772 42140
rect 16604 42084 16660 42094
rect 16604 41990 16660 42028
rect 16716 41746 16772 41758
rect 16716 41694 16718 41746
rect 16770 41694 16772 41746
rect 16380 41188 16436 41198
rect 16156 40740 16212 40750
rect 16156 40514 16212 40684
rect 16380 40626 16436 41132
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 16380 40562 16436 40574
rect 16156 40462 16158 40514
rect 16210 40462 16212 40514
rect 16156 40450 16212 40462
rect 16604 40404 16660 40414
rect 16492 40402 16660 40404
rect 16492 40350 16606 40402
rect 16658 40350 16660 40402
rect 16492 40348 16660 40350
rect 16492 40292 16548 40348
rect 16604 40338 16660 40348
rect 16380 39618 16436 39630
rect 16380 39566 16382 39618
rect 16434 39566 16436 39618
rect 16380 39508 16436 39566
rect 16380 39442 16436 39452
rect 16492 39396 16548 40236
rect 16716 39844 16772 41694
rect 16492 39330 16548 39340
rect 16604 39788 16772 39844
rect 17164 41186 17220 41198
rect 17164 41134 17166 41186
rect 17218 41134 17220 41186
rect 15820 37490 15988 37492
rect 15820 37438 15822 37490
rect 15874 37438 15988 37490
rect 15820 37436 15988 37438
rect 16044 38164 16100 38174
rect 15820 37426 15876 37436
rect 16044 37380 16100 38108
rect 16156 37940 16212 37950
rect 16156 37604 16212 37884
rect 16380 37826 16436 37838
rect 16380 37774 16382 37826
rect 16434 37774 16436 37826
rect 16380 37604 16436 37774
rect 16492 37604 16548 37614
rect 16380 37548 16492 37604
rect 16156 37538 16212 37548
rect 16492 37538 16548 37548
rect 16044 37314 16100 37324
rect 16268 37378 16324 37390
rect 16268 37326 16270 37378
rect 16322 37326 16324 37378
rect 15932 37268 15988 37278
rect 15932 37174 15988 37212
rect 16156 37268 16212 37278
rect 16268 37268 16324 37326
rect 16492 37380 16548 37390
rect 16492 37286 16548 37324
rect 16212 37212 16324 37268
rect 16156 37202 16212 37212
rect 15708 37100 15876 37156
rect 15820 37044 15876 37100
rect 16156 37044 16212 37054
rect 15820 36988 16100 37044
rect 15484 36754 15540 36764
rect 15036 35870 15038 35922
rect 15090 35870 15092 35922
rect 15036 35858 15092 35870
rect 15260 35812 15316 35822
rect 15148 35588 15204 35598
rect 15260 35588 15316 35756
rect 15204 35532 15316 35588
rect 15372 35588 15428 35598
rect 15148 35522 15204 35532
rect 14812 35026 14980 35028
rect 14812 34974 14814 35026
rect 14866 34974 14980 35026
rect 14812 34972 14980 34974
rect 14812 34962 14868 34972
rect 14364 34402 14420 34412
rect 14476 34412 14644 34468
rect 14700 34914 14756 34926
rect 14700 34862 14702 34914
rect 14754 34862 14756 34914
rect 14364 34242 14420 34254
rect 14364 34190 14366 34242
rect 14418 34190 14420 34242
rect 14364 33124 14420 34190
rect 14364 33058 14420 33068
rect 14364 32676 14420 32686
rect 14364 32582 14420 32620
rect 14476 31948 14532 34412
rect 14700 34020 14756 34862
rect 14924 34804 14980 34814
rect 14924 34710 14980 34748
rect 15148 34804 15204 34814
rect 15036 34580 15092 34590
rect 14700 33954 14756 33964
rect 14812 34468 14868 34478
rect 14812 34242 14868 34412
rect 14812 34190 14814 34242
rect 14866 34190 14868 34242
rect 14588 33124 14644 33134
rect 14588 33030 14644 33068
rect 14812 33012 14868 34190
rect 15036 33570 15092 34524
rect 15036 33518 15038 33570
rect 15090 33518 15092 33570
rect 15036 33458 15092 33518
rect 15036 33406 15038 33458
rect 15090 33406 15092 33458
rect 15036 33394 15092 33406
rect 15148 34468 15204 34748
rect 15260 34468 15316 34478
rect 15148 34412 15260 34468
rect 15148 33236 15204 34412
rect 15260 34402 15316 34412
rect 15260 34132 15316 34142
rect 15260 34038 15316 34076
rect 15148 33180 15316 33236
rect 14812 32956 15092 33012
rect 14924 32788 14980 32798
rect 14812 32452 14868 32462
rect 14252 31154 14308 31164
rect 14364 31892 14532 31948
rect 14700 32450 14868 32452
rect 14700 32398 14814 32450
rect 14866 32398 14868 32450
rect 14700 32396 14868 32398
rect 14364 31218 14420 31892
rect 14588 31668 14644 31678
rect 14364 31166 14366 31218
rect 14418 31166 14420 31218
rect 14252 30882 14308 30894
rect 14252 30830 14254 30882
rect 14306 30830 14308 30882
rect 14028 30716 14196 30772
rect 13804 29810 13860 29820
rect 14028 30210 14084 30222
rect 14028 30158 14030 30210
rect 14082 30158 14084 30210
rect 14028 30100 14084 30158
rect 14140 30100 14196 30716
rect 14252 30212 14308 30830
rect 14364 30434 14420 31166
rect 14364 30382 14366 30434
rect 14418 30382 14420 30434
rect 14364 30370 14420 30382
rect 14476 31666 14644 31668
rect 14476 31614 14590 31666
rect 14642 31614 14644 31666
rect 14476 31612 14644 31614
rect 14476 30324 14532 31612
rect 14588 31602 14644 31612
rect 14588 30996 14644 31006
rect 14700 30996 14756 32396
rect 14812 32386 14868 32396
rect 14924 32004 14980 32732
rect 15036 32340 15092 32956
rect 15036 32274 15092 32284
rect 14924 31938 14980 31948
rect 15148 32004 15204 32014
rect 14812 31668 14868 31678
rect 14812 31574 14868 31612
rect 15036 31668 15092 31678
rect 15148 31668 15204 31948
rect 15260 31778 15316 33180
rect 15260 31726 15262 31778
rect 15314 31726 15316 31778
rect 15260 31714 15316 31726
rect 15036 31666 15204 31668
rect 15036 31614 15038 31666
rect 15090 31614 15204 31666
rect 15036 31612 15204 31614
rect 15036 31602 15092 31612
rect 14924 31556 14980 31566
rect 14924 31462 14980 31500
rect 14588 30994 14756 30996
rect 14588 30942 14590 30994
rect 14642 30942 14756 30994
rect 14588 30940 14756 30942
rect 14588 30930 14644 30940
rect 14700 30772 14756 30940
rect 14700 30706 14756 30716
rect 14812 31332 14868 31342
rect 14812 30660 14868 31276
rect 15148 31220 15204 31230
rect 15148 31126 15204 31164
rect 14812 30594 14868 30604
rect 15148 30770 15204 30782
rect 15148 30718 15150 30770
rect 15202 30718 15204 30770
rect 14924 30434 14980 30446
rect 14924 30382 14926 30434
rect 14978 30382 14980 30434
rect 14476 30268 14868 30324
rect 14252 30156 14756 30212
rect 14140 30044 14308 30100
rect 13692 29540 13748 29550
rect 13244 29372 13524 29428
rect 13132 29362 13188 29372
rect 13020 28030 13022 28082
rect 13074 28030 13076 28082
rect 13020 28018 13076 28030
rect 13132 29202 13188 29214
rect 13132 29150 13134 29202
rect 13186 29150 13188 29202
rect 13132 28084 13188 29150
rect 13356 29202 13412 29214
rect 13356 29150 13358 29202
rect 13410 29150 13412 29202
rect 13356 28756 13412 29150
rect 13356 28690 13412 28700
rect 13468 28532 13524 29372
rect 13692 29092 13748 29484
rect 13916 29428 13972 29438
rect 13804 29372 13916 29428
rect 13804 29202 13860 29372
rect 13916 29362 13972 29372
rect 13804 29150 13806 29202
rect 13858 29150 13860 29202
rect 13804 29138 13860 29150
rect 13916 29204 13972 29214
rect 14028 29204 14084 30044
rect 13916 29202 14084 29204
rect 13916 29150 13918 29202
rect 13970 29150 14084 29202
rect 13916 29148 14084 29150
rect 13916 29138 13972 29148
rect 13692 29026 13748 29036
rect 13132 28018 13188 28028
rect 13356 28476 13524 28532
rect 13356 26908 13412 28476
rect 14140 28196 14196 28206
rect 13692 28084 13748 28094
rect 13692 27858 13748 28028
rect 13692 27806 13694 27858
rect 13746 27806 13748 27858
rect 13692 27794 13748 27806
rect 14028 27858 14084 27870
rect 14028 27806 14030 27858
rect 14082 27806 14084 27858
rect 14028 27748 14084 27806
rect 12908 26852 13076 26908
rect 12796 26674 12852 26684
rect 12796 26516 12852 26526
rect 12796 25508 12852 26460
rect 12908 25508 12964 25518
rect 12796 25506 12964 25508
rect 12796 25454 12910 25506
rect 12962 25454 12964 25506
rect 12796 25452 12964 25454
rect 12908 25442 12964 25452
rect 12572 25396 12628 25406
rect 12572 25302 12628 25340
rect 12796 25282 12852 25294
rect 12796 25230 12798 25282
rect 12850 25230 12852 25282
rect 12796 24948 12852 25230
rect 13020 25172 13076 26852
rect 13244 26852 13412 26908
rect 13580 26964 13636 27002
rect 14028 26908 14084 27692
rect 14140 27186 14196 28140
rect 14140 27134 14142 27186
rect 14194 27134 14196 27186
rect 14140 27122 14196 27134
rect 13580 26898 13636 26908
rect 13804 26852 14084 26908
rect 13244 26516 13300 26852
rect 13244 26422 13300 26460
rect 13692 26516 13748 26526
rect 13692 26422 13748 26460
rect 13580 26292 13636 26302
rect 13356 25172 13412 25182
rect 13020 25116 13188 25172
rect 13020 24948 13076 24958
rect 12796 24892 13020 24948
rect 13020 24722 13076 24892
rect 13020 24670 13022 24722
rect 13074 24670 13076 24722
rect 13020 24658 13076 24670
rect 13132 24724 13188 25116
rect 13132 24500 13188 24668
rect 12460 23998 12462 24050
rect 12514 23998 12516 24050
rect 12460 23828 12516 23998
rect 12908 24444 13188 24500
rect 13356 24722 13412 25116
rect 13356 24670 13358 24722
rect 13410 24670 13412 24722
rect 12908 23938 12964 24444
rect 12908 23886 12910 23938
rect 12962 23886 12964 23938
rect 12908 23874 12964 23886
rect 12460 23762 12516 23772
rect 11340 23538 11396 23548
rect 13356 23492 13412 24670
rect 13580 24722 13636 26236
rect 13692 25284 13748 25294
rect 13692 25190 13748 25228
rect 13804 25172 13860 26852
rect 14252 26628 14308 30044
rect 14476 29986 14532 29998
rect 14476 29934 14478 29986
rect 14530 29934 14532 29986
rect 14364 29876 14420 29886
rect 14476 29876 14532 29934
rect 14420 29820 14532 29876
rect 14364 29810 14420 29820
rect 14700 29538 14756 30156
rect 14700 29486 14702 29538
rect 14754 29486 14756 29538
rect 14700 29474 14756 29486
rect 14812 29652 14868 30268
rect 14924 30322 14980 30382
rect 14924 30270 14926 30322
rect 14978 30270 14980 30322
rect 14924 29764 14980 30270
rect 14924 29698 14980 29708
rect 14364 29428 14420 29438
rect 14364 29334 14420 29372
rect 14588 29426 14644 29438
rect 14588 29374 14590 29426
rect 14642 29374 14644 29426
rect 14476 28980 14532 28990
rect 14588 28980 14644 29374
rect 14812 29428 14868 29596
rect 15148 29650 15204 30718
rect 15148 29598 15150 29650
rect 15202 29598 15204 29650
rect 15148 29586 15204 29598
rect 15372 29428 15428 35532
rect 15820 34802 15876 34814
rect 15820 34750 15822 34802
rect 15874 34750 15876 34802
rect 15820 34354 15876 34750
rect 15820 34302 15822 34354
rect 15874 34302 15876 34354
rect 15820 34290 15876 34302
rect 15484 34244 15540 34254
rect 15484 33458 15540 34188
rect 15932 34242 15988 34254
rect 15932 34190 15934 34242
rect 15986 34190 15988 34242
rect 15484 33406 15486 33458
rect 15538 33406 15540 33458
rect 15484 33394 15540 33406
rect 15820 34132 15876 34142
rect 15484 32452 15540 32462
rect 15484 32358 15540 32396
rect 15708 32452 15764 32462
rect 15484 31780 15540 31790
rect 15484 31218 15540 31724
rect 15484 31166 15486 31218
rect 15538 31166 15540 31218
rect 15484 30884 15540 31166
rect 15484 30818 15540 30828
rect 15708 30770 15764 32396
rect 15820 32004 15876 34076
rect 15932 33908 15988 34190
rect 16044 34132 16100 36988
rect 16156 36950 16212 36988
rect 16380 37044 16436 37054
rect 16156 34132 16212 34142
rect 16044 34130 16212 34132
rect 16044 34078 16158 34130
rect 16210 34078 16212 34130
rect 16044 34076 16212 34078
rect 15932 33012 15988 33852
rect 15932 32946 15988 32956
rect 16156 33236 16212 34076
rect 16380 33348 16436 36988
rect 16604 37044 16660 39788
rect 16940 37938 16996 37950
rect 16940 37886 16942 37938
rect 16994 37886 16996 37938
rect 16828 37828 16884 37838
rect 16940 37828 16996 37886
rect 16884 37772 16996 37828
rect 16828 37762 16884 37772
rect 16604 36978 16660 36988
rect 16828 37492 16884 37502
rect 16604 36372 16660 36382
rect 16492 34914 16548 34926
rect 16492 34862 16494 34914
rect 16546 34862 16548 34914
rect 16492 33460 16548 34862
rect 16604 34244 16660 36316
rect 16828 35308 16884 37436
rect 17164 37492 17220 41134
rect 17500 40402 17556 43148
rect 18060 42980 18116 43708
rect 18172 43428 18228 47292
rect 18284 47124 18340 47406
rect 18396 47460 18452 47470
rect 18396 47366 18452 47404
rect 18508 47124 18564 48524
rect 18620 47684 18676 48748
rect 18844 48738 18900 48748
rect 19180 48354 19236 49086
rect 19964 49138 20020 49150
rect 19964 49086 19966 49138
rect 20018 49086 20020 49138
rect 19180 48302 19182 48354
rect 19234 48302 19236 48354
rect 19180 48290 19236 48302
rect 19404 49026 19460 49038
rect 19404 48974 19406 49026
rect 19458 48974 19460 49026
rect 19404 48020 19460 48974
rect 19964 49028 20020 49086
rect 19964 48962 20020 48972
rect 20524 49026 20580 49196
rect 20524 48974 20526 49026
rect 20578 48974 20580 49026
rect 20524 48962 20580 48974
rect 19628 48916 19684 48926
rect 19628 48822 19684 48860
rect 19852 48914 19908 48926
rect 19852 48862 19854 48914
rect 19906 48862 19908 48914
rect 19740 48804 19796 48814
rect 19852 48804 19908 48862
rect 20412 48916 20468 48926
rect 20412 48822 20468 48860
rect 19796 48748 19908 48804
rect 20188 48802 20244 48814
rect 20188 48750 20190 48802
rect 20242 48750 20244 48802
rect 19740 48738 19796 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19964 48466 20020 48478
rect 20188 48468 20244 48750
rect 19964 48414 19966 48466
rect 20018 48414 20020 48466
rect 19852 48354 19908 48366
rect 19852 48302 19854 48354
rect 19906 48302 19908 48354
rect 19852 48132 19908 48302
rect 19852 48066 19908 48076
rect 19404 47954 19460 47964
rect 18620 47682 19460 47684
rect 18620 47630 18622 47682
rect 18674 47630 19460 47682
rect 18620 47628 19460 47630
rect 18620 47618 18676 47628
rect 19180 47460 19236 47470
rect 19180 47366 19236 47404
rect 19404 47460 19460 47628
rect 19404 47404 19908 47460
rect 18284 47068 18564 47124
rect 18396 44324 18452 44334
rect 18396 44230 18452 44268
rect 18508 43708 18564 47068
rect 18732 47346 18788 47358
rect 18732 47294 18734 47346
rect 18786 47294 18788 47346
rect 18620 44994 18676 45006
rect 18620 44942 18622 44994
rect 18674 44942 18676 44994
rect 18620 44884 18676 44942
rect 18620 43876 18676 44828
rect 18620 43810 18676 43820
rect 18284 43652 18340 43662
rect 18396 43652 18564 43708
rect 18340 43596 18452 43652
rect 18620 43650 18676 43662
rect 18620 43598 18622 43650
rect 18674 43598 18676 43650
rect 18284 43586 18340 43596
rect 18508 43540 18564 43550
rect 18508 43446 18564 43484
rect 18172 43372 18340 43428
rect 17612 42924 18116 42980
rect 17612 42754 17668 42924
rect 17612 42702 17614 42754
rect 17666 42702 17668 42754
rect 17612 42196 17668 42702
rect 17612 42130 17668 42140
rect 17836 42756 17892 42766
rect 17836 42082 17892 42700
rect 18060 42754 18116 42766
rect 18060 42702 18062 42754
rect 18114 42702 18116 42754
rect 18060 42532 18116 42702
rect 18060 42308 18116 42476
rect 18060 42242 18116 42252
rect 17836 42030 17838 42082
rect 17890 42030 17892 42082
rect 17836 42018 17892 42030
rect 17948 42084 18004 42094
rect 17948 41972 18004 42028
rect 18284 41972 18340 43372
rect 18620 42420 18676 43598
rect 18620 42354 18676 42364
rect 18508 42084 18564 42094
rect 17948 41916 18116 41972
rect 17836 41860 17892 41870
rect 17836 41748 17892 41804
rect 17948 41748 18004 41758
rect 17836 41746 18004 41748
rect 17836 41694 17950 41746
rect 18002 41694 18004 41746
rect 17836 41692 18004 41694
rect 17948 41682 18004 41692
rect 18060 41524 18116 41916
rect 17948 41468 18116 41524
rect 18172 41916 18340 41972
rect 18396 41970 18452 41982
rect 18396 41918 18398 41970
rect 18450 41918 18452 41970
rect 17612 41188 17668 41198
rect 17612 41094 17668 41132
rect 17500 40350 17502 40402
rect 17554 40350 17556 40402
rect 17500 40180 17556 40350
rect 17500 40114 17556 40124
rect 17724 40514 17780 40526
rect 17724 40462 17726 40514
rect 17778 40462 17780 40514
rect 17724 40180 17780 40462
rect 17724 40114 17780 40124
rect 17836 40516 17892 40526
rect 17388 39732 17444 39742
rect 17388 39618 17444 39676
rect 17388 39566 17390 39618
rect 17442 39566 17444 39618
rect 17388 39554 17444 39566
rect 17836 39284 17892 40460
rect 17836 39218 17892 39228
rect 17948 38276 18004 41468
rect 18172 41298 18228 41916
rect 18396 41860 18452 41918
rect 18172 41246 18174 41298
rect 18226 41246 18228 41298
rect 18172 41234 18228 41246
rect 18284 41804 18452 41860
rect 18172 40852 18228 40862
rect 18172 40626 18228 40796
rect 18172 40574 18174 40626
rect 18226 40574 18228 40626
rect 18172 40562 18228 40574
rect 18060 40516 18116 40526
rect 18060 39394 18116 40460
rect 18060 39342 18062 39394
rect 18114 39342 18116 39394
rect 18060 39330 18116 39342
rect 18172 39506 18228 39518
rect 18172 39454 18174 39506
rect 18226 39454 18228 39506
rect 18172 39060 18228 39454
rect 18172 38994 18228 39004
rect 18060 38724 18116 38734
rect 18284 38668 18340 41804
rect 18508 41748 18564 42028
rect 18620 41972 18676 41982
rect 18732 41972 18788 47294
rect 19404 47346 19460 47404
rect 19404 47294 19406 47346
rect 19458 47294 19460 47346
rect 19404 47282 19460 47294
rect 19852 47346 19908 47404
rect 19852 47294 19854 47346
rect 19906 47294 19908 47346
rect 19852 47282 19908 47294
rect 19292 47234 19348 47246
rect 19740 47236 19796 47246
rect 19292 47182 19294 47234
rect 19346 47182 19348 47234
rect 19292 46676 19348 47182
rect 19292 46610 19348 46620
rect 19516 47234 19796 47236
rect 19516 47182 19742 47234
rect 19794 47182 19796 47234
rect 19516 47180 19796 47182
rect 19964 47236 20020 48414
rect 20076 48412 20244 48468
rect 20076 48242 20132 48412
rect 20076 48190 20078 48242
rect 20130 48190 20132 48242
rect 20076 48178 20132 48190
rect 20524 48132 20580 48142
rect 20300 48020 20356 48030
rect 20076 47460 20132 47470
rect 20076 47366 20132 47404
rect 20300 47460 20356 47964
rect 20300 47366 20356 47404
rect 19964 47180 20244 47236
rect 19516 46004 19572 47180
rect 19740 47170 19796 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 46900 20244 47180
rect 20524 47124 20580 48076
rect 20524 47058 20580 47068
rect 20076 46844 20244 46900
rect 20076 46116 20132 46844
rect 20748 46786 20804 46798
rect 20748 46734 20750 46786
rect 20802 46734 20804 46786
rect 20748 46452 20804 46734
rect 20076 46060 20244 46116
rect 19180 45948 19572 46004
rect 18844 45892 18900 45902
rect 18844 42084 18900 45836
rect 18844 42018 18900 42028
rect 18956 45220 19012 45230
rect 18620 41970 18788 41972
rect 18620 41918 18622 41970
rect 18674 41918 18788 41970
rect 18620 41916 18788 41918
rect 18956 41972 19012 45164
rect 19068 45218 19124 45230
rect 19068 45166 19070 45218
rect 19122 45166 19124 45218
rect 19068 44996 19124 45166
rect 19068 44322 19124 44940
rect 19068 44270 19070 44322
rect 19122 44270 19124 44322
rect 19068 43764 19124 44270
rect 19068 43698 19124 43708
rect 18956 41916 19124 41972
rect 18620 41906 18676 41916
rect 18844 41858 18900 41870
rect 18844 41806 18846 41858
rect 18898 41806 18900 41858
rect 18508 41692 18788 41748
rect 18620 40852 18676 40862
rect 18620 40514 18676 40796
rect 18620 40462 18622 40514
rect 18674 40462 18676 40514
rect 18620 40450 18676 40462
rect 18508 40292 18564 40302
rect 18732 40292 18788 41692
rect 18844 41412 18900 41806
rect 18844 41346 18900 41356
rect 18956 41746 19012 41758
rect 18956 41694 18958 41746
rect 19010 41694 19012 41746
rect 18508 40198 18564 40236
rect 18620 40236 18788 40292
rect 18844 40402 18900 40414
rect 18844 40350 18846 40402
rect 18898 40350 18900 40402
rect 18060 38630 18116 38668
rect 18172 38612 18340 38668
rect 18396 38612 18452 38622
rect 17948 38220 18116 38276
rect 17164 37426 17220 37436
rect 17276 38050 17332 38062
rect 17276 37998 17278 38050
rect 17330 37998 17332 38050
rect 17276 37268 17332 37998
rect 17948 38052 18004 38062
rect 17948 37958 18004 37996
rect 17836 37940 17892 37950
rect 17836 37846 17892 37884
rect 17164 36820 17220 36830
rect 16828 35252 17108 35308
rect 16828 35140 16884 35150
rect 16828 34802 16884 35084
rect 17052 35026 17108 35252
rect 17052 34974 17054 35026
rect 17106 34974 17108 35026
rect 17052 34962 17108 34974
rect 16940 34916 16996 34926
rect 16940 34822 16996 34860
rect 16828 34750 16830 34802
rect 16882 34750 16884 34802
rect 16828 34738 16884 34750
rect 16604 34178 16660 34188
rect 16716 34132 16772 34142
rect 16716 34038 16772 34076
rect 17052 33460 17108 33470
rect 16492 33404 16660 33460
rect 16156 33012 16212 33180
rect 16156 32946 16212 32956
rect 16268 33292 16436 33348
rect 15820 31948 15988 32004
rect 15820 31780 15876 31790
rect 15820 31686 15876 31724
rect 15708 30718 15710 30770
rect 15762 30718 15764 30770
rect 15708 30706 15764 30718
rect 15484 30660 15540 30670
rect 15484 30210 15540 30604
rect 15484 30158 15486 30210
rect 15538 30158 15540 30210
rect 15484 30146 15540 30158
rect 15932 29764 15988 31948
rect 16044 31666 16100 31678
rect 16044 31614 16046 31666
rect 16098 31614 16100 31666
rect 16044 31108 16100 31614
rect 16268 31220 16324 33292
rect 16380 33122 16436 33134
rect 16380 33070 16382 33122
rect 16434 33070 16436 33122
rect 16380 33012 16436 33070
rect 16380 32946 16436 32956
rect 16604 32676 16660 33404
rect 17052 33236 17108 33404
rect 17164 33458 17220 36764
rect 17276 34354 17332 37212
rect 17388 37826 17444 37838
rect 17388 37774 17390 37826
rect 17442 37774 17444 37826
rect 17388 37156 17444 37774
rect 17612 37828 17668 37838
rect 17948 37828 18004 37838
rect 17612 37826 17780 37828
rect 17612 37774 17614 37826
rect 17666 37774 17780 37826
rect 17612 37772 17780 37774
rect 17612 37762 17668 37772
rect 17388 37090 17444 37100
rect 17500 37604 17556 37614
rect 17500 37268 17556 37548
rect 17612 37268 17668 37278
rect 17556 37266 17668 37268
rect 17556 37214 17614 37266
rect 17666 37214 17668 37266
rect 17556 37212 17668 37214
rect 17500 36594 17556 37212
rect 17612 37202 17668 37212
rect 17500 36542 17502 36594
rect 17554 36542 17556 36594
rect 17500 36530 17556 36542
rect 17724 36036 17780 37772
rect 17948 37716 18004 37772
rect 17836 37660 18004 37716
rect 17836 36484 17892 37660
rect 17948 37492 18004 37502
rect 18060 37492 18116 38220
rect 17948 37490 18116 37492
rect 17948 37438 17950 37490
rect 18002 37438 18116 37490
rect 17948 37436 18116 37438
rect 17948 37426 18004 37436
rect 18060 36708 18116 37436
rect 18060 36642 18116 36652
rect 18172 36706 18228 38612
rect 18396 38050 18452 38556
rect 18396 37998 18398 38050
rect 18450 37998 18452 38050
rect 18396 37986 18452 37998
rect 18508 38052 18564 38062
rect 18508 37958 18564 37996
rect 18620 37604 18676 40236
rect 18732 39620 18788 39630
rect 18732 39526 18788 39564
rect 18844 39060 18900 40350
rect 18956 40404 19012 41694
rect 18956 40338 19012 40348
rect 18732 39004 18900 39060
rect 18732 38276 18788 39004
rect 19068 38948 19124 41916
rect 19180 39172 19236 45948
rect 19964 45892 20020 45902
rect 19404 45890 20020 45892
rect 19404 45838 19966 45890
rect 20018 45838 20020 45890
rect 19404 45836 20020 45838
rect 19404 45218 19460 45836
rect 19964 45826 20020 45836
rect 20076 45892 20132 45902
rect 20076 45798 20132 45836
rect 19740 45668 19796 45678
rect 19628 45666 19796 45668
rect 19628 45614 19742 45666
rect 19794 45614 19796 45666
rect 19628 45612 19796 45614
rect 19404 45166 19406 45218
rect 19458 45166 19460 45218
rect 19292 44212 19348 44222
rect 19404 44212 19460 45166
rect 19516 45220 19572 45230
rect 19628 45220 19684 45612
rect 19740 45602 19796 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19572 45164 19684 45220
rect 19740 45330 19796 45342
rect 20188 45332 20244 46060
rect 19740 45278 19742 45330
rect 19794 45278 19796 45330
rect 19516 45154 19572 45164
rect 19740 44996 19796 45278
rect 20076 45276 20244 45332
rect 20636 45666 20692 45678
rect 20636 45614 20638 45666
rect 20690 45614 20692 45666
rect 19292 44210 19460 44212
rect 19292 44158 19294 44210
rect 19346 44158 19460 44210
rect 19292 44156 19460 44158
rect 19628 44940 19796 44996
rect 19964 45106 20020 45118
rect 19964 45054 19966 45106
rect 20018 45054 20020 45106
rect 19292 44146 19348 44156
rect 19628 43652 19684 44940
rect 19964 44772 20020 45054
rect 19964 44706 20020 44716
rect 20076 44100 20132 45276
rect 20636 45220 20692 45614
rect 20748 45444 20804 46396
rect 21308 46674 21364 46686
rect 21308 46622 21310 46674
rect 21362 46622 21364 46674
rect 20748 45378 20804 45388
rect 20860 46004 20916 46014
rect 20412 45164 20692 45220
rect 20748 45220 20804 45230
rect 20300 44996 20356 45006
rect 20412 44996 20468 45164
rect 20748 45106 20804 45164
rect 20748 45054 20750 45106
rect 20802 45054 20804 45106
rect 20748 45042 20804 45054
rect 20300 44994 20468 44996
rect 20300 44942 20302 44994
rect 20354 44942 20468 44994
rect 20300 44940 20468 44942
rect 20524 44996 20580 45006
rect 20300 44212 20356 44940
rect 20524 44902 20580 44940
rect 20300 44146 20356 44156
rect 20076 44044 20244 44100
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19628 43586 19684 43596
rect 20188 43540 20244 44044
rect 20524 43540 20580 43550
rect 20188 43538 20580 43540
rect 20188 43486 20526 43538
rect 20578 43486 20580 43538
rect 20188 43484 20580 43486
rect 20524 43474 20580 43484
rect 20412 42868 20468 42878
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19404 42196 19460 42206
rect 19404 41074 19460 42140
rect 19964 42084 20020 42094
rect 19964 41970 20020 42028
rect 19964 41918 19966 41970
rect 20018 41918 20020 41970
rect 19964 41906 20020 41918
rect 20300 41970 20356 41982
rect 20300 41918 20302 41970
rect 20354 41918 20356 41970
rect 19852 41860 19908 41870
rect 19404 41022 19406 41074
rect 19458 41022 19460 41074
rect 19404 41010 19460 41022
rect 19516 41636 19572 41646
rect 19516 40626 19572 41580
rect 19628 41412 19684 41422
rect 19628 41186 19684 41356
rect 19628 41134 19630 41186
rect 19682 41134 19684 41186
rect 19628 41122 19684 41134
rect 19852 41188 19908 41804
rect 20300 41860 20356 41918
rect 20300 41794 20356 41804
rect 19964 41188 20020 41198
rect 19852 41186 20020 41188
rect 19852 41134 19966 41186
rect 20018 41134 20020 41186
rect 19852 41132 20020 41134
rect 19964 41122 20020 41132
rect 19852 40964 19908 41002
rect 19852 40898 19908 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19516 40574 19518 40626
rect 19570 40574 19572 40626
rect 19516 40562 19572 40574
rect 19292 40404 19348 40442
rect 19292 40338 19348 40348
rect 19628 40404 19684 40414
rect 19180 39106 19236 39116
rect 19292 40180 19348 40190
rect 19068 38892 19236 38948
rect 18844 38724 18900 38734
rect 18844 38500 18900 38668
rect 19180 38668 19236 38892
rect 19292 38836 19348 40124
rect 19628 39956 19684 40348
rect 19516 39900 19684 39956
rect 19404 39844 19460 39854
rect 19404 39284 19460 39788
rect 19404 39058 19460 39228
rect 19404 39006 19406 39058
rect 19458 39006 19460 39058
rect 19404 38994 19460 39006
rect 19292 38770 19348 38780
rect 19180 38612 19460 38668
rect 18844 38444 19236 38500
rect 19068 38276 19124 38286
rect 18732 38274 19124 38276
rect 18732 38222 19070 38274
rect 19122 38222 19124 38274
rect 18732 38220 19124 38222
rect 19068 38210 19124 38220
rect 18508 37548 18676 37604
rect 18732 38050 18788 38062
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18284 37492 18340 37502
rect 18284 37378 18340 37436
rect 18284 37326 18286 37378
rect 18338 37326 18340 37378
rect 18284 37314 18340 37326
rect 18396 37378 18452 37390
rect 18396 37326 18398 37378
rect 18450 37326 18452 37378
rect 18396 36932 18452 37326
rect 18396 36866 18452 36876
rect 18172 36654 18174 36706
rect 18226 36654 18228 36706
rect 18172 36642 18228 36654
rect 18060 36484 18116 36494
rect 17836 36428 18004 36484
rect 17836 36260 17892 36270
rect 17836 36166 17892 36204
rect 17724 35980 17892 36036
rect 17724 35810 17780 35822
rect 17724 35758 17726 35810
rect 17778 35758 17780 35810
rect 17612 35700 17668 35710
rect 17276 34302 17278 34354
rect 17330 34302 17332 34354
rect 17276 34290 17332 34302
rect 17388 35698 17668 35700
rect 17388 35646 17614 35698
rect 17666 35646 17668 35698
rect 17388 35644 17668 35646
rect 17164 33406 17166 33458
rect 17218 33406 17220 33458
rect 17164 33394 17220 33406
rect 17276 33572 17332 33582
rect 17052 33170 17108 33180
rect 17164 33234 17220 33246
rect 17164 33182 17166 33234
rect 17218 33182 17220 33234
rect 17164 33124 17220 33182
rect 16268 31126 16324 31164
rect 16380 32620 16660 32676
rect 16828 32676 16884 32686
rect 16044 30884 16100 31052
rect 16044 30818 16100 30828
rect 16156 30994 16212 31006
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 16156 30212 16212 30942
rect 16268 30884 16324 30894
rect 16268 30770 16324 30828
rect 16268 30718 16270 30770
rect 16322 30718 16324 30770
rect 16268 30706 16324 30718
rect 16156 29988 16212 30156
rect 16156 29922 16212 29932
rect 15932 29708 16212 29764
rect 15708 29652 15764 29662
rect 15764 29596 16100 29652
rect 15708 29558 15764 29596
rect 15372 29372 15988 29428
rect 14812 29362 14868 29372
rect 15372 29204 15428 29214
rect 15148 29202 15428 29204
rect 15148 29150 15374 29202
rect 15426 29150 15428 29202
rect 15148 29148 15428 29150
rect 14588 28924 14756 28980
rect 14476 28754 14532 28924
rect 14700 28868 14756 28924
rect 14700 28812 15092 28868
rect 14476 28702 14478 28754
rect 14530 28702 14532 28754
rect 14476 28690 14532 28702
rect 15036 28754 15092 28812
rect 15036 28702 15038 28754
rect 15090 28702 15092 28754
rect 15036 28690 15092 28702
rect 15148 28642 15204 29148
rect 15372 29138 15428 29148
rect 15148 28590 15150 28642
rect 15202 28590 15204 28642
rect 14700 28530 14756 28542
rect 14700 28478 14702 28530
rect 14754 28478 14756 28530
rect 14700 28084 14756 28478
rect 14924 28420 14980 28430
rect 14924 28326 14980 28364
rect 15148 28308 15204 28590
rect 15260 28980 15316 28990
rect 15260 28642 15316 28924
rect 15260 28590 15262 28642
rect 15314 28590 15316 28642
rect 15260 28578 15316 28590
rect 15148 28242 15204 28252
rect 14364 27412 14420 27422
rect 14364 26964 14420 27356
rect 14476 27076 14532 27086
rect 14476 26982 14532 27020
rect 14700 27074 14756 28028
rect 15484 27860 15540 27870
rect 15708 27860 15764 27870
rect 15484 27766 15540 27804
rect 15596 27858 15764 27860
rect 15596 27806 15710 27858
rect 15762 27806 15764 27858
rect 15596 27804 15764 27806
rect 14924 27412 14980 27422
rect 15596 27412 15652 27804
rect 15708 27794 15764 27804
rect 15820 27858 15876 27870
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15820 27636 15876 27806
rect 15820 27570 15876 27580
rect 14700 27022 14702 27074
rect 14754 27022 14756 27074
rect 14700 27010 14756 27022
rect 14812 27356 14924 27412
rect 14364 26898 14420 26908
rect 14140 26516 14196 26526
rect 14252 26516 14308 26572
rect 14140 26514 14308 26516
rect 14140 26462 14142 26514
rect 14194 26462 14308 26514
rect 14140 26460 14308 26462
rect 14140 26450 14196 26460
rect 14028 25508 14084 25518
rect 14028 25394 14084 25452
rect 14252 25506 14308 26460
rect 14700 26516 14756 26526
rect 14812 26516 14868 27356
rect 14924 27346 14980 27356
rect 15260 27356 15652 27412
rect 15708 27412 15764 27422
rect 15260 27186 15316 27356
rect 15260 27134 15262 27186
rect 15314 27134 15316 27186
rect 15260 27122 15316 27134
rect 14924 27076 14980 27086
rect 14924 26908 14980 27020
rect 15148 27076 15204 27086
rect 15148 26982 15204 27020
rect 15708 27074 15764 27356
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15708 27010 15764 27022
rect 15372 26964 15428 27002
rect 14924 26852 15092 26908
rect 15372 26898 15428 26908
rect 15820 26962 15876 26974
rect 15820 26910 15822 26962
rect 15874 26910 15876 26962
rect 15036 26796 15204 26852
rect 14700 26514 14868 26516
rect 14700 26462 14702 26514
rect 14754 26462 14868 26514
rect 14700 26460 14868 26462
rect 14700 26450 14756 26460
rect 15036 26404 15092 26414
rect 15036 26310 15092 26348
rect 14924 25620 14980 25630
rect 14924 25526 14980 25564
rect 14252 25454 14254 25506
rect 14306 25454 14308 25506
rect 14252 25442 14308 25454
rect 14028 25342 14030 25394
rect 14082 25342 14084 25394
rect 14028 25330 14084 25342
rect 13804 25106 13860 25116
rect 14028 25060 14084 25070
rect 13580 24670 13582 24722
rect 13634 24670 13636 24722
rect 13580 24658 13636 24670
rect 13916 24724 13972 24734
rect 13916 24630 13972 24668
rect 14028 24050 14084 25004
rect 14028 23998 14030 24050
rect 14082 23998 14084 24050
rect 14028 23986 14084 23998
rect 14700 24948 14756 24958
rect 14700 23938 14756 24892
rect 15148 24836 15204 26796
rect 15596 26740 15652 26750
rect 15484 26516 15540 26526
rect 15484 26290 15540 26460
rect 15596 26514 15652 26684
rect 15596 26462 15598 26514
rect 15650 26462 15652 26514
rect 15596 26450 15652 26462
rect 15708 26404 15764 26414
rect 15708 26310 15764 26348
rect 15484 26238 15486 26290
rect 15538 26238 15540 26290
rect 15484 26226 15540 26238
rect 15820 26290 15876 26910
rect 15820 26238 15822 26290
rect 15874 26238 15876 26290
rect 15260 25620 15316 25630
rect 15260 25506 15316 25564
rect 15820 25620 15876 26238
rect 15932 26740 15988 29372
rect 16044 28642 16100 29596
rect 16156 29650 16212 29708
rect 16156 29598 16158 29650
rect 16210 29598 16212 29650
rect 16156 29202 16212 29598
rect 16156 29150 16158 29202
rect 16210 29150 16212 29202
rect 16156 29138 16212 29150
rect 16044 28590 16046 28642
rect 16098 28590 16100 28642
rect 16044 28578 16100 28590
rect 16268 28084 16324 28094
rect 16268 27990 16324 28028
rect 16380 27300 16436 32620
rect 16828 32582 16884 32620
rect 16492 32450 16548 32462
rect 16492 32398 16494 32450
rect 16546 32398 16548 32450
rect 16492 32004 16548 32398
rect 16492 31938 16548 31948
rect 16604 31778 16660 31790
rect 16604 31726 16606 31778
rect 16658 31726 16660 31778
rect 16604 31444 16660 31726
rect 17052 31778 17108 31790
rect 17052 31726 17054 31778
rect 17106 31726 17108 31778
rect 17052 31668 17108 31726
rect 16604 31378 16660 31388
rect 16716 31612 17108 31668
rect 16716 29316 16772 31612
rect 16044 27244 16436 27300
rect 16492 29260 16772 29316
rect 16828 30882 16884 30894
rect 16828 30830 16830 30882
rect 16882 30830 16884 30882
rect 16828 30660 16884 30830
rect 16044 27074 16100 27244
rect 16044 27022 16046 27074
rect 16098 27022 16100 27074
rect 16044 27010 16100 27022
rect 15932 26068 15988 26684
rect 16492 26404 16548 29260
rect 16604 29092 16660 29102
rect 16604 28754 16660 29036
rect 16604 28702 16606 28754
rect 16658 28702 16660 28754
rect 16604 28420 16660 28702
rect 16604 28354 16660 28364
rect 16716 28308 16772 28318
rect 16716 28082 16772 28252
rect 16716 28030 16718 28082
rect 16770 28030 16772 28082
rect 16716 28018 16772 28030
rect 16604 27858 16660 27870
rect 16604 27806 16606 27858
rect 16658 27806 16660 27858
rect 16604 27412 16660 27806
rect 16716 27636 16772 27646
rect 16716 27542 16772 27580
rect 16828 27524 16884 30604
rect 17052 30100 17108 30110
rect 17164 30100 17220 33068
rect 17276 31108 17332 33516
rect 17388 32002 17444 35644
rect 17612 35634 17668 35644
rect 17724 35476 17780 35758
rect 17724 35410 17780 35420
rect 17724 35252 17780 35262
rect 17500 34244 17556 34254
rect 17500 34150 17556 34188
rect 17612 34130 17668 34142
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17612 34020 17668 34078
rect 17388 31950 17390 32002
rect 17442 31950 17444 32002
rect 17388 31938 17444 31950
rect 17500 33964 17612 34020
rect 17388 31108 17444 31118
rect 17276 31106 17444 31108
rect 17276 31054 17390 31106
rect 17442 31054 17444 31106
rect 17276 31052 17444 31054
rect 17388 31042 17444 31052
rect 17276 30548 17332 30558
rect 17276 30210 17332 30492
rect 17276 30158 17278 30210
rect 17330 30158 17332 30210
rect 17276 30146 17332 30158
rect 17500 30210 17556 33964
rect 17612 33954 17668 33964
rect 17612 33460 17668 33470
rect 17612 33346 17668 33404
rect 17612 33294 17614 33346
rect 17666 33294 17668 33346
rect 17612 33282 17668 33294
rect 17612 32900 17668 32910
rect 17724 32900 17780 35196
rect 17836 35028 17892 35980
rect 17836 34962 17892 34972
rect 17836 34692 17892 34702
rect 17836 33348 17892 34636
rect 17948 33572 18004 36428
rect 18060 36390 18116 36428
rect 18284 36370 18340 36382
rect 18284 36318 18286 36370
rect 18338 36318 18340 36370
rect 18284 34804 18340 36318
rect 18396 35924 18452 35934
rect 18396 35588 18452 35868
rect 18396 35522 18452 35532
rect 18284 34738 18340 34748
rect 18508 35140 18564 37548
rect 18620 37268 18676 37278
rect 18732 37268 18788 37998
rect 18620 37266 18788 37268
rect 18620 37214 18622 37266
rect 18674 37214 18788 37266
rect 18620 37212 18788 37214
rect 18844 38052 18900 38062
rect 18620 37202 18676 37212
rect 18508 34692 18564 35084
rect 18508 34626 18564 34636
rect 18620 36708 18676 36718
rect 18060 34580 18116 34590
rect 18060 34354 18116 34524
rect 18060 34302 18062 34354
rect 18114 34302 18116 34354
rect 18060 34132 18116 34302
rect 18508 34356 18564 34366
rect 18620 34356 18676 36652
rect 18732 36706 18788 36718
rect 18732 36654 18734 36706
rect 18786 36654 18788 36706
rect 18732 35922 18788 36654
rect 18844 36596 18900 37996
rect 18956 38050 19012 38062
rect 18956 37998 18958 38050
rect 19010 37998 19012 38050
rect 18956 37828 19012 37998
rect 18956 37762 19012 37772
rect 19068 37940 19124 37950
rect 18844 36502 18900 36540
rect 18956 37380 19012 37390
rect 18956 36372 19012 37324
rect 18732 35870 18734 35922
rect 18786 35870 18788 35922
rect 18732 35858 18788 35870
rect 18844 36316 19012 36372
rect 19068 37266 19124 37884
rect 19068 37214 19070 37266
rect 19122 37214 19124 37266
rect 18732 35698 18788 35710
rect 18732 35646 18734 35698
rect 18786 35646 18788 35698
rect 18732 35026 18788 35646
rect 18844 35252 18900 36316
rect 19068 35588 19124 37214
rect 19180 37378 19236 38444
rect 19180 37326 19182 37378
rect 19234 37326 19236 37378
rect 19180 36932 19236 37326
rect 19180 36866 19236 36876
rect 19292 38052 19348 38062
rect 19180 35812 19236 35822
rect 19180 35718 19236 35756
rect 19292 35700 19348 37996
rect 19404 37604 19460 38612
rect 19404 37538 19460 37548
rect 19404 37380 19460 37390
rect 19516 37380 19572 39900
rect 20412 39620 20468 42812
rect 20748 42084 20804 42094
rect 20748 41990 20804 42028
rect 20524 41970 20580 41982
rect 20524 41918 20526 41970
rect 20578 41918 20580 41970
rect 20524 41074 20580 41918
rect 20860 41972 20916 45948
rect 21308 45332 21364 46622
rect 21420 45892 21476 50372
rect 22428 50034 22484 50372
rect 22764 50260 22820 50372
rect 22764 50194 22820 50204
rect 22428 49982 22430 50034
rect 22482 49982 22484 50034
rect 22428 49970 22484 49982
rect 22204 49924 22260 49934
rect 22092 49810 22148 49822
rect 22092 49758 22094 49810
rect 22146 49758 22148 49810
rect 21756 49700 21812 49710
rect 22092 49700 22148 49758
rect 21812 49644 22148 49700
rect 21756 49606 21812 49644
rect 21532 49252 21588 49262
rect 21532 48356 21588 49196
rect 21868 49028 21924 49038
rect 21868 48934 21924 48972
rect 22092 49026 22148 49038
rect 22092 48974 22094 49026
rect 22146 48974 22148 49026
rect 21532 48354 21700 48356
rect 21532 48302 21534 48354
rect 21586 48302 21700 48354
rect 21532 48300 21700 48302
rect 21532 48290 21588 48300
rect 21420 45826 21476 45836
rect 21532 47460 21588 47470
rect 21532 46674 21588 47404
rect 21644 47012 21700 48300
rect 21868 48354 21924 48366
rect 21868 48302 21870 48354
rect 21922 48302 21924 48354
rect 21868 48020 21924 48302
rect 22092 48244 22148 48974
rect 22204 49026 22260 49868
rect 23324 49588 23380 55356
rect 25452 55300 25508 55310
rect 25564 55300 25620 56142
rect 25788 56082 25844 56364
rect 25788 56030 25790 56082
rect 25842 56030 25844 56082
rect 25788 56018 25844 56030
rect 27580 55858 27636 59200
rect 29820 56420 29876 59200
rect 29820 56364 30324 56420
rect 29820 56306 29876 56364
rect 29820 56254 29822 56306
rect 29874 56254 29876 56306
rect 29820 56242 29876 56254
rect 28364 56196 28420 56206
rect 27580 55806 27582 55858
rect 27634 55806 27636 55858
rect 27580 55794 27636 55806
rect 27692 56194 28420 56196
rect 27692 56142 28366 56194
rect 28418 56142 28420 56194
rect 27692 56140 28420 56142
rect 25452 55298 25620 55300
rect 25452 55246 25454 55298
rect 25506 55246 25620 55298
rect 25452 55244 25620 55246
rect 27692 55298 27748 56140
rect 28364 56130 28420 56140
rect 30044 56194 30100 56206
rect 30044 56142 30046 56194
rect 30098 56142 30100 56194
rect 28588 56082 28644 56094
rect 28588 56030 28590 56082
rect 28642 56030 28644 56082
rect 27916 55972 27972 55982
rect 27916 55858 27972 55916
rect 28588 55972 28644 56030
rect 28588 55906 28644 55916
rect 27916 55806 27918 55858
rect 27970 55806 27972 55858
rect 27916 55794 27972 55806
rect 28364 55860 28420 55870
rect 27692 55246 27694 55298
rect 27746 55246 27748 55298
rect 25452 55234 25508 55244
rect 27692 55234 27748 55246
rect 25340 55074 25396 55086
rect 25340 55022 25342 55074
rect 25394 55022 25396 55074
rect 23436 54516 23492 54526
rect 23436 53170 23492 54460
rect 25228 54514 25284 54526
rect 25228 54462 25230 54514
rect 25282 54462 25284 54514
rect 23884 54402 23940 54414
rect 23884 54350 23886 54402
rect 23938 54350 23940 54402
rect 23660 53844 23716 53854
rect 23660 53750 23716 53788
rect 23436 53118 23438 53170
rect 23490 53118 23492 53170
rect 23436 53106 23492 53118
rect 23548 53506 23604 53518
rect 23548 53454 23550 53506
rect 23602 53454 23604 53506
rect 23548 52052 23604 53454
rect 23548 51986 23604 51996
rect 23772 53508 23828 53518
rect 23884 53508 23940 54350
rect 24780 54404 24836 54414
rect 24444 53730 24500 53742
rect 24444 53678 24446 53730
rect 24498 53678 24500 53730
rect 23772 53506 23940 53508
rect 23772 53454 23774 53506
rect 23826 53454 23940 53506
rect 23772 53452 23940 53454
rect 23996 53506 24052 53518
rect 23996 53454 23998 53506
rect 24050 53454 24052 53506
rect 22204 48974 22206 49026
rect 22258 48974 22260 49026
rect 22204 48962 22260 48974
rect 22988 49532 23380 49588
rect 23548 51492 23604 51502
rect 22540 48914 22596 48926
rect 22876 48916 22932 48926
rect 22540 48862 22542 48914
rect 22594 48862 22596 48914
rect 22428 48802 22484 48814
rect 22428 48750 22430 48802
rect 22482 48750 22484 48802
rect 22428 48356 22484 48750
rect 22428 48290 22484 48300
rect 22092 48178 22148 48188
rect 22316 48244 22372 48254
rect 22316 48132 22372 48188
rect 22428 48132 22484 48142
rect 22316 48130 22484 48132
rect 22316 48078 22430 48130
rect 22482 48078 22484 48130
rect 22316 48076 22484 48078
rect 22204 48020 22260 48030
rect 21868 48018 22260 48020
rect 21868 47966 22206 48018
rect 22258 47966 22260 48018
rect 21868 47964 22260 47966
rect 21644 46946 21700 46956
rect 21532 46622 21534 46674
rect 21586 46622 21588 46674
rect 21532 45890 21588 46622
rect 22092 46676 22148 46686
rect 22092 46582 22148 46620
rect 21532 45838 21534 45890
rect 21586 45838 21588 45890
rect 21420 45332 21476 45342
rect 21308 45330 21476 45332
rect 21308 45278 21422 45330
rect 21474 45278 21476 45330
rect 21308 45276 21476 45278
rect 21532 45332 21588 45838
rect 21868 46340 21924 46350
rect 21756 45780 21812 45790
rect 21756 45686 21812 45724
rect 21644 45332 21700 45342
rect 21532 45330 21700 45332
rect 21532 45278 21646 45330
rect 21698 45278 21700 45330
rect 21532 45276 21700 45278
rect 21420 45266 21476 45276
rect 21644 45266 21700 45276
rect 20972 44884 21028 44894
rect 20972 44790 21028 44828
rect 21420 44324 21476 44334
rect 21420 44098 21476 44268
rect 21420 44046 21422 44098
rect 21474 44046 21476 44098
rect 21420 43988 21476 44046
rect 21420 43922 21476 43932
rect 21868 44212 21924 46284
rect 22204 46002 22260 47964
rect 22316 46228 22372 48076
rect 22428 48066 22484 48076
rect 22540 48020 22596 48862
rect 22764 48914 22932 48916
rect 22764 48862 22878 48914
rect 22930 48862 22932 48914
rect 22764 48860 22932 48862
rect 22764 48242 22820 48860
rect 22876 48850 22932 48860
rect 22988 48914 23044 49532
rect 22988 48862 22990 48914
rect 23042 48862 23044 48914
rect 22988 48850 23044 48862
rect 23212 48802 23268 48814
rect 23212 48750 23214 48802
rect 23266 48750 23268 48802
rect 23212 48468 23268 48750
rect 23212 48402 23268 48412
rect 22764 48190 22766 48242
rect 22818 48190 22820 48242
rect 22764 48020 22820 48190
rect 22540 48018 22820 48020
rect 22540 47966 22542 48018
rect 22594 47966 22820 48018
rect 22540 47964 22820 47966
rect 22876 48354 22932 48366
rect 22876 48302 22878 48354
rect 22930 48302 22932 48354
rect 22540 47954 22596 47964
rect 22876 47236 22932 48302
rect 22876 47170 22932 47180
rect 22988 48356 23044 48366
rect 22652 47012 22708 47022
rect 22652 46786 22708 46956
rect 22652 46734 22654 46786
rect 22706 46734 22708 46786
rect 22652 46722 22708 46734
rect 22316 46162 22372 46172
rect 22428 46562 22484 46574
rect 22428 46510 22430 46562
rect 22482 46510 22484 46562
rect 22428 46004 22484 46510
rect 22204 45950 22206 46002
rect 22258 45950 22260 46002
rect 22204 45938 22260 45950
rect 22316 45948 22484 46004
rect 20972 43876 21028 43886
rect 20972 42194 21028 43820
rect 21644 43652 21700 43662
rect 21644 43650 21812 43652
rect 21644 43598 21646 43650
rect 21698 43598 21812 43650
rect 21644 43596 21812 43598
rect 21644 43586 21700 43596
rect 21756 43540 21812 43596
rect 21756 43474 21812 43484
rect 21756 42868 21812 42878
rect 21308 42532 21364 42542
rect 21308 42438 21364 42476
rect 20972 42142 20974 42194
rect 21026 42142 21028 42194
rect 20972 42130 21028 42142
rect 20972 41972 21028 41982
rect 20860 41970 21028 41972
rect 20860 41918 20974 41970
rect 21026 41918 21028 41970
rect 20860 41916 21028 41918
rect 20972 41860 21028 41916
rect 20972 41794 21028 41804
rect 21532 41858 21588 41870
rect 21532 41806 21534 41858
rect 21586 41806 21588 41858
rect 21532 41748 21588 41806
rect 21532 41682 21588 41692
rect 21756 41636 21812 42812
rect 21868 41748 21924 44156
rect 21980 45890 22036 45902
rect 21980 45838 21982 45890
rect 22034 45838 22036 45890
rect 21980 43876 22036 45838
rect 22092 45892 22148 45902
rect 22092 45332 22148 45836
rect 22316 45444 22372 45948
rect 22428 45780 22484 45790
rect 22428 45686 22484 45724
rect 22540 45668 22596 45678
rect 22540 45666 22820 45668
rect 22540 45614 22542 45666
rect 22594 45614 22820 45666
rect 22540 45612 22820 45614
rect 22540 45602 22596 45612
rect 22316 45388 22484 45444
rect 22092 45276 22372 45332
rect 22316 45218 22372 45276
rect 22316 45166 22318 45218
rect 22370 45166 22372 45218
rect 22316 45154 22372 45166
rect 22092 45106 22148 45118
rect 22092 45054 22094 45106
rect 22146 45054 22148 45106
rect 22092 44772 22148 45054
rect 22092 44706 22148 44716
rect 22204 45106 22260 45118
rect 22204 45054 22206 45106
rect 22258 45054 22260 45106
rect 22204 44436 22260 45054
rect 22204 44370 22260 44380
rect 21980 43810 22036 43820
rect 22092 43988 22148 43998
rect 22092 43540 22148 43932
rect 22204 43764 22260 43774
rect 22204 43670 22260 43708
rect 22092 43484 22372 43540
rect 21980 41972 22036 41982
rect 21980 41878 22036 41916
rect 22092 41970 22148 41982
rect 22092 41918 22094 41970
rect 22146 41918 22148 41970
rect 21868 41692 22036 41748
rect 21756 41580 21924 41636
rect 21756 41412 21812 41422
rect 21308 41410 21812 41412
rect 21308 41358 21758 41410
rect 21810 41358 21812 41410
rect 21308 41356 21812 41358
rect 20860 41188 20916 41198
rect 21308 41188 21364 41356
rect 21756 41346 21812 41356
rect 20860 41186 21364 41188
rect 20860 41134 20862 41186
rect 20914 41134 21364 41186
rect 20860 41132 21364 41134
rect 21420 41188 21476 41226
rect 20860 41122 20916 41132
rect 21420 41122 21476 41132
rect 21532 41186 21588 41198
rect 21532 41134 21534 41186
rect 21586 41134 21588 41186
rect 20524 41022 20526 41074
rect 20578 41022 20580 41074
rect 20524 40964 20580 41022
rect 20524 40898 20580 40908
rect 20636 40962 20692 40974
rect 20636 40910 20638 40962
rect 20690 40910 20692 40962
rect 20636 40180 20692 40910
rect 21084 40964 21140 40974
rect 21084 40626 21140 40908
rect 21084 40574 21086 40626
rect 21138 40574 21140 40626
rect 21084 40562 21140 40574
rect 21532 40404 21588 41134
rect 21532 40338 21588 40348
rect 20692 40124 21028 40180
rect 20636 40114 20692 40124
rect 20412 39554 20468 39564
rect 19628 39508 19684 39518
rect 19628 39414 19684 39452
rect 20300 39396 20356 39406
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19964 38722 20020 38734
rect 19964 38670 19966 38722
rect 20018 38670 20020 38722
rect 19964 38668 20020 38670
rect 19740 38612 19796 38622
rect 19628 38556 19740 38612
rect 19628 38162 19684 38556
rect 19740 38546 19796 38556
rect 19852 38612 20020 38668
rect 20300 38722 20356 39340
rect 20972 38834 21028 40124
rect 21308 39620 21364 39630
rect 21308 39526 21364 39564
rect 20972 38782 20974 38834
rect 21026 38782 21028 38834
rect 20972 38770 21028 38782
rect 21084 39060 21140 39070
rect 20300 38670 20302 38722
rect 20354 38670 20356 38722
rect 20300 38612 20356 38670
rect 21084 38668 21140 39004
rect 21196 39004 21812 39060
rect 21196 38834 21252 39004
rect 21196 38782 21198 38834
rect 21250 38782 21252 38834
rect 21196 38770 21252 38782
rect 21308 38834 21364 38846
rect 21308 38782 21310 38834
rect 21362 38782 21364 38834
rect 21308 38668 21364 38782
rect 21532 38834 21588 38846
rect 21532 38782 21534 38834
rect 21586 38782 21588 38834
rect 21532 38668 21588 38782
rect 21756 38668 21812 39004
rect 21084 38612 21364 38668
rect 21420 38612 21588 38668
rect 21644 38612 21812 38668
rect 19628 38110 19630 38162
rect 19682 38110 19684 38162
rect 19628 38098 19684 38110
rect 19740 38164 19796 38174
rect 19852 38164 19908 38612
rect 19796 38108 19908 38164
rect 19740 38098 19796 38108
rect 19964 38052 20020 38062
rect 19964 37958 20020 37996
rect 19740 37940 19796 37950
rect 19740 37846 19796 37884
rect 20188 37940 20244 37950
rect 19404 37378 19572 37380
rect 19404 37326 19406 37378
rect 19458 37326 19572 37378
rect 19404 37324 19572 37326
rect 19628 37828 19684 37838
rect 19404 37314 19460 37324
rect 19404 37156 19460 37166
rect 19460 37100 19572 37156
rect 19404 37090 19460 37100
rect 19404 36258 19460 36270
rect 19404 36206 19406 36258
rect 19458 36206 19460 36258
rect 19404 36036 19460 36206
rect 19404 35970 19460 35980
rect 19516 35812 19572 37100
rect 19628 35924 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 37884
rect 20076 37436 20244 37492
rect 20076 37380 20132 37436
rect 20076 37314 20132 37324
rect 20076 37156 20132 37166
rect 20076 36706 20132 37100
rect 20300 37044 20356 38556
rect 21420 38388 21476 38612
rect 20636 38332 21476 38388
rect 20636 38274 20692 38332
rect 20636 38222 20638 38274
rect 20690 38222 20692 38274
rect 20636 38210 20692 38222
rect 20300 36978 20356 36988
rect 20412 38050 20468 38062
rect 20412 37998 20414 38050
rect 20466 37998 20468 38050
rect 20076 36654 20078 36706
rect 20130 36654 20132 36706
rect 20076 36642 20132 36654
rect 20412 36482 20468 37998
rect 21420 37828 21476 37838
rect 21308 37826 21476 37828
rect 21308 37774 21422 37826
rect 21474 37774 21476 37826
rect 21308 37772 21476 37774
rect 20860 37716 20916 37726
rect 20860 37266 20916 37660
rect 20860 37214 20862 37266
rect 20914 37214 20916 37266
rect 20860 37202 20916 37214
rect 21084 37268 21140 37278
rect 21308 37268 21364 37772
rect 21420 37762 21476 37772
rect 21644 37492 21700 38612
rect 21084 37266 21364 37268
rect 21084 37214 21086 37266
rect 21138 37214 21364 37266
rect 21084 37212 21364 37214
rect 21420 37436 21700 37492
rect 21868 37826 21924 41580
rect 21980 41410 22036 41692
rect 21980 41358 21982 41410
rect 22034 41358 22036 41410
rect 21980 40964 22036 41358
rect 22092 41410 22148 41918
rect 22204 41970 22260 41982
rect 22204 41918 22206 41970
rect 22258 41918 22260 41970
rect 22204 41748 22260 41918
rect 22204 41682 22260 41692
rect 22092 41358 22094 41410
rect 22146 41358 22148 41410
rect 22092 41346 22148 41358
rect 21980 40898 22036 40908
rect 22204 39620 22260 39630
rect 21980 39060 22036 39070
rect 21980 38966 22036 39004
rect 22204 39058 22260 39564
rect 22204 39006 22206 39058
rect 22258 39006 22260 39058
rect 22204 38994 22260 39006
rect 21868 37774 21870 37826
rect 21922 37774 21924 37826
rect 21084 37044 21140 37212
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 20412 36418 20468 36430
rect 20748 36988 21140 37044
rect 20748 36596 20804 36988
rect 20748 36482 20804 36540
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20748 36418 20804 36430
rect 20860 36484 20916 36494
rect 20188 36372 20244 36382
rect 19740 36260 19796 36298
rect 20188 36278 20244 36316
rect 19740 36194 19796 36204
rect 20412 36260 20468 36270
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35924 19796 35934
rect 19628 35922 19796 35924
rect 19628 35870 19742 35922
rect 19794 35870 19796 35922
rect 19628 35868 19796 35870
rect 19740 35858 19796 35868
rect 19516 35756 19684 35812
rect 19292 35644 19572 35700
rect 19068 35532 19236 35588
rect 18844 35196 19012 35252
rect 18732 34974 18734 35026
rect 18786 34974 18788 35026
rect 18732 34962 18788 34974
rect 18844 34804 18900 34814
rect 18844 34710 18900 34748
rect 18956 34580 19012 35196
rect 19068 34692 19124 34730
rect 19068 34626 19124 34636
rect 18844 34524 19012 34580
rect 18620 34300 18788 34356
rect 18508 34262 18564 34300
rect 18396 34132 18452 34142
rect 18060 34066 18116 34076
rect 18284 34130 18452 34132
rect 18284 34078 18398 34130
rect 18450 34078 18452 34130
rect 18284 34076 18452 34078
rect 18284 33908 18340 34076
rect 18396 34066 18452 34076
rect 18620 34130 18676 34142
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 17948 33506 18004 33516
rect 18060 33852 18340 33908
rect 17836 33292 18004 33348
rect 17668 32844 17780 32900
rect 17836 32900 17892 32910
rect 17612 32834 17668 32844
rect 17724 32676 17780 32686
rect 17724 32562 17780 32620
rect 17724 32510 17726 32562
rect 17778 32510 17780 32562
rect 17724 32498 17780 32510
rect 17836 32116 17892 32844
rect 17948 32674 18004 33292
rect 17948 32622 17950 32674
rect 18002 32622 18004 32674
rect 17948 32610 18004 32622
rect 17836 32050 17892 32060
rect 17948 32340 18004 32350
rect 18060 32340 18116 33852
rect 18508 33346 18564 33358
rect 18508 33294 18510 33346
rect 18562 33294 18564 33346
rect 18284 33122 18340 33134
rect 18284 33070 18286 33122
rect 18338 33070 18340 33122
rect 18284 32900 18340 33070
rect 18284 32834 18340 32844
rect 18004 32284 18116 32340
rect 18172 32450 18228 32462
rect 18172 32398 18174 32450
rect 18226 32398 18228 32450
rect 17724 31778 17780 31790
rect 17724 31726 17726 31778
rect 17778 31726 17780 31778
rect 17612 31108 17668 31118
rect 17612 31014 17668 31052
rect 17500 30158 17502 30210
rect 17554 30158 17556 30210
rect 17108 30044 17220 30100
rect 17052 30034 17108 30044
rect 17500 29092 17556 30158
rect 17724 30884 17780 31726
rect 17948 31666 18004 32284
rect 18172 32004 18228 32398
rect 18172 31938 18228 31948
rect 18284 31892 18340 31902
rect 18284 31798 18340 31836
rect 18508 31780 18564 33294
rect 18620 33124 18676 34078
rect 18620 33058 18676 33068
rect 18508 31686 18564 31724
rect 18620 32340 18676 32350
rect 17948 31614 17950 31666
rect 18002 31614 18004 31666
rect 17948 31602 18004 31614
rect 17836 31556 17892 31566
rect 17836 31218 17892 31500
rect 18060 31556 18116 31566
rect 17836 31166 17838 31218
rect 17890 31166 17892 31218
rect 17836 31154 17892 31166
rect 17948 31444 18004 31454
rect 17724 29876 17780 30828
rect 17500 29026 17556 29036
rect 17612 29820 17780 29876
rect 17836 30996 17892 31006
rect 17500 28868 17556 28878
rect 16828 27458 16884 27468
rect 17052 28420 17108 28430
rect 17052 27412 17108 28364
rect 16604 27356 16772 27412
rect 16492 26338 16548 26348
rect 16604 26850 16660 26862
rect 16604 26798 16606 26850
rect 16658 26798 16660 26850
rect 16044 26292 16100 26302
rect 16044 26198 16100 26236
rect 16156 26180 16212 26190
rect 16604 26180 16660 26798
rect 16212 26124 16324 26180
rect 16156 26114 16212 26124
rect 15932 26002 15988 26012
rect 15820 25554 15876 25564
rect 15260 25454 15262 25506
rect 15314 25454 15316 25506
rect 15260 25442 15316 25454
rect 16044 25508 16100 25518
rect 16044 25414 16100 25452
rect 15260 25284 15316 25294
rect 15260 25190 15316 25228
rect 16044 24836 16100 24846
rect 15148 24834 16100 24836
rect 15148 24782 16046 24834
rect 16098 24782 16100 24834
rect 15148 24780 16100 24782
rect 15596 24276 15652 24286
rect 15148 24052 15204 24062
rect 15148 23958 15204 23996
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14700 23874 14756 23886
rect 15596 23938 15652 24220
rect 15596 23886 15598 23938
rect 15650 23886 15652 23938
rect 13356 23426 13412 23436
rect 15148 23828 15204 23838
rect 15148 23378 15204 23772
rect 15148 23326 15150 23378
rect 15202 23326 15204 23378
rect 15148 23314 15204 23326
rect 15596 23378 15652 23886
rect 15596 23326 15598 23378
rect 15650 23326 15652 23378
rect 15596 23314 15652 23326
rect 15932 23828 15988 23838
rect 15932 23378 15988 23772
rect 15932 23326 15934 23378
rect 15986 23326 15988 23378
rect 15932 23314 15988 23326
rect 8316 23202 8372 23212
rect 15820 23268 15876 23278
rect 15820 23174 15876 23212
rect 16044 22932 16100 24780
rect 16156 24052 16212 24062
rect 16268 24052 16324 26124
rect 16604 26114 16660 26124
rect 16380 25620 16436 25630
rect 16380 25394 16436 25564
rect 16492 25620 16548 25630
rect 16492 25618 16660 25620
rect 16492 25566 16494 25618
rect 16546 25566 16660 25618
rect 16492 25564 16660 25566
rect 16492 25554 16548 25564
rect 16380 25342 16382 25394
rect 16434 25342 16436 25394
rect 16380 25330 16436 25342
rect 16492 24722 16548 24734
rect 16492 24670 16494 24722
rect 16546 24670 16548 24722
rect 16492 24612 16548 24670
rect 16492 24546 16548 24556
rect 16156 24050 16324 24052
rect 16156 23998 16158 24050
rect 16210 23998 16324 24050
rect 16156 23996 16324 23998
rect 16156 23986 16212 23996
rect 16380 23938 16436 23950
rect 16380 23886 16382 23938
rect 16434 23886 16436 23938
rect 16380 23492 16436 23886
rect 16156 23436 16436 23492
rect 16492 23828 16548 23838
rect 16604 23828 16660 25564
rect 16716 25508 16772 27356
rect 17052 27346 17108 27356
rect 17164 28308 17220 28318
rect 17164 27186 17220 28252
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 16716 25442 16772 25452
rect 16828 26178 16884 26190
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 25396 16884 26126
rect 16716 24946 16772 24958
rect 16716 24894 16718 24946
rect 16770 24894 16772 24946
rect 16716 24724 16772 24894
rect 16716 24658 16772 24668
rect 16828 24612 16884 25340
rect 16940 26068 16996 26078
rect 16940 24836 16996 26012
rect 16940 24770 16996 24780
rect 17164 24836 17220 27134
rect 17388 27524 17444 27534
rect 17388 26908 17444 27468
rect 17500 27076 17556 28812
rect 17612 27298 17668 29820
rect 17612 27246 17614 27298
rect 17666 27246 17668 27298
rect 17612 27234 17668 27246
rect 17724 27858 17780 27870
rect 17724 27806 17726 27858
rect 17778 27806 17780 27858
rect 17500 27010 17556 27020
rect 17612 26962 17668 26974
rect 17612 26910 17614 26962
rect 17666 26910 17668 26962
rect 17612 26908 17668 26910
rect 17388 26852 17668 26908
rect 17612 26740 17668 26750
rect 17612 26404 17668 26684
rect 17724 26514 17780 27806
rect 17836 27634 17892 30940
rect 17948 30548 18004 31388
rect 18060 31106 18116 31500
rect 18060 31054 18062 31106
rect 18114 31054 18116 31106
rect 18060 31042 18116 31054
rect 18620 30994 18676 32284
rect 18732 31220 18788 34300
rect 18844 32900 18900 34524
rect 19068 34468 19124 34478
rect 19068 34130 19124 34412
rect 19068 34078 19070 34130
rect 19122 34078 19124 34130
rect 19068 34018 19124 34078
rect 19068 33966 19070 34018
rect 19122 33966 19124 34018
rect 19068 33954 19124 33966
rect 18956 33572 19012 33582
rect 19180 33572 19236 35532
rect 19292 35028 19348 35038
rect 19292 34914 19348 34972
rect 19292 34862 19294 34914
rect 19346 34862 19348 34914
rect 19292 34850 19348 34862
rect 19404 34914 19460 34926
rect 19404 34862 19406 34914
rect 19458 34862 19460 34914
rect 18956 33570 19236 33572
rect 18956 33518 18958 33570
rect 19010 33518 19236 33570
rect 18956 33516 19236 33518
rect 19292 34020 19348 34030
rect 18956 33506 19012 33516
rect 19292 33460 19348 33964
rect 19068 33234 19124 33246
rect 19068 33182 19070 33234
rect 19122 33182 19124 33234
rect 18956 33124 19012 33134
rect 18956 33030 19012 33068
rect 18844 32844 19012 32900
rect 18844 32564 18900 32574
rect 18844 32470 18900 32508
rect 18956 32340 19012 32844
rect 19068 32564 19124 33182
rect 19180 32788 19236 32798
rect 19292 32788 19348 33404
rect 19180 32786 19348 32788
rect 19180 32734 19182 32786
rect 19234 32734 19348 32786
rect 19180 32732 19348 32734
rect 19180 32722 19236 32732
rect 19068 32498 19124 32508
rect 18956 32284 19236 32340
rect 18956 31668 19012 31678
rect 18956 31554 19012 31612
rect 18956 31502 18958 31554
rect 19010 31502 19012 31554
rect 18956 31444 19012 31502
rect 18956 31378 19012 31388
rect 19068 31220 19124 31230
rect 18732 31218 19124 31220
rect 18732 31166 19070 31218
rect 19122 31166 19124 31218
rect 18732 31164 19124 31166
rect 19068 31108 19124 31164
rect 19068 31042 19124 31052
rect 18620 30942 18622 30994
rect 18674 30942 18676 30994
rect 18620 30930 18676 30942
rect 18732 30994 18788 31006
rect 18732 30942 18734 30994
rect 18786 30942 18788 30994
rect 18172 30884 18228 30894
rect 18172 30790 18228 30828
rect 17948 30482 18004 30492
rect 18284 30212 18340 30222
rect 18284 30118 18340 30156
rect 18732 30212 18788 30942
rect 18956 30994 19012 31006
rect 18956 30942 18958 30994
rect 19010 30942 19012 30994
rect 18844 30884 18900 30894
rect 18844 30790 18900 30828
rect 18956 30660 19012 30942
rect 19180 30884 19236 32284
rect 18956 30594 19012 30604
rect 19068 30828 19236 30884
rect 18732 30146 18788 30156
rect 18956 29652 19012 29662
rect 18732 29596 18956 29652
rect 18620 29540 18676 29550
rect 18508 28644 18564 28654
rect 18172 28642 18564 28644
rect 18172 28590 18510 28642
rect 18562 28590 18564 28642
rect 18172 28588 18564 28590
rect 18172 28082 18228 28588
rect 18508 28578 18564 28588
rect 18284 28420 18340 28430
rect 18620 28420 18676 29484
rect 18284 28326 18340 28364
rect 18396 28364 18676 28420
rect 18732 29316 18788 29596
rect 18956 29558 19012 29596
rect 18732 28530 18788 29260
rect 18844 28644 18900 28654
rect 18844 28550 18900 28588
rect 18732 28478 18734 28530
rect 18786 28478 18788 28530
rect 18732 28420 18788 28478
rect 18172 28030 18174 28082
rect 18226 28030 18228 28082
rect 18172 28018 18228 28030
rect 18396 27970 18452 28364
rect 18732 28354 18788 28364
rect 18396 27918 18398 27970
rect 18450 27918 18452 27970
rect 18396 27906 18452 27918
rect 17948 27860 18004 27870
rect 17948 27858 18340 27860
rect 17948 27806 17950 27858
rect 18002 27806 18340 27858
rect 17948 27804 18340 27806
rect 17948 27794 18004 27804
rect 17836 27582 17838 27634
rect 17890 27582 17892 27634
rect 17836 27570 17892 27582
rect 18060 27412 18116 27422
rect 17724 26462 17726 26514
rect 17778 26462 17780 26514
rect 17724 26450 17780 26462
rect 17836 27298 17892 27310
rect 17836 27246 17838 27298
rect 17890 27246 17892 27298
rect 17612 26310 17668 26348
rect 17388 26290 17444 26302
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 17388 26180 17444 26238
rect 17388 25506 17444 26124
rect 17836 26290 17892 27246
rect 17948 27300 18004 27310
rect 17948 26516 18004 27244
rect 18060 27188 18116 27356
rect 18284 27188 18340 27804
rect 18732 27858 18788 27870
rect 18732 27806 18734 27858
rect 18786 27806 18788 27858
rect 18620 27524 18676 27534
rect 18508 27188 18564 27198
rect 18284 27186 18564 27188
rect 18284 27134 18510 27186
rect 18562 27134 18564 27186
rect 18284 27132 18564 27134
rect 18060 27094 18116 27132
rect 18508 27122 18564 27132
rect 18620 27074 18676 27468
rect 18732 27412 18788 27806
rect 18732 27346 18788 27356
rect 18620 27022 18622 27074
rect 18674 27022 18676 27074
rect 18620 27010 18676 27022
rect 18844 27076 18900 27086
rect 18396 26964 18452 27002
rect 18396 26898 18452 26908
rect 18844 26962 18900 27020
rect 18844 26910 18846 26962
rect 18898 26910 18900 26962
rect 18844 26898 18900 26910
rect 19068 26908 19124 30828
rect 19292 30660 19348 30670
rect 19292 30210 19348 30604
rect 19404 30324 19460 34862
rect 19516 34692 19572 35644
rect 19516 34626 19572 34636
rect 19628 34132 19684 35756
rect 19964 35810 20020 35822
rect 19964 35758 19966 35810
rect 20018 35758 20020 35810
rect 19852 35588 19908 35598
rect 19852 34916 19908 35532
rect 19964 35476 20020 35758
rect 20076 35700 20132 35710
rect 20076 35698 20244 35700
rect 20076 35646 20078 35698
rect 20130 35646 20244 35698
rect 20076 35644 20244 35646
rect 20076 35634 20132 35644
rect 19964 35420 20132 35476
rect 20076 35308 20132 35420
rect 19852 34850 19908 34860
rect 19964 35252 20132 35308
rect 19964 34692 20020 35252
rect 20188 35140 20244 35644
rect 20076 35084 20244 35140
rect 20300 35252 20356 35262
rect 20076 34916 20132 35084
rect 20076 34850 20132 34860
rect 20188 34916 20244 34926
rect 20300 34916 20356 35196
rect 20188 34914 20356 34916
rect 20188 34862 20190 34914
rect 20242 34862 20356 34914
rect 20188 34860 20356 34862
rect 20412 34914 20468 36204
rect 20636 36258 20692 36270
rect 20636 36206 20638 36258
rect 20690 36206 20692 36258
rect 20412 34862 20414 34914
rect 20466 34862 20468 34914
rect 20188 34850 20244 34860
rect 20412 34850 20468 34862
rect 20524 35810 20580 35822
rect 20524 35758 20526 35810
rect 20578 35758 20580 35810
rect 20300 34692 20356 34702
rect 19964 34690 20356 34692
rect 19964 34638 20302 34690
rect 20354 34638 20356 34690
rect 19964 34636 20356 34638
rect 20300 34626 20356 34636
rect 20412 34580 20468 34590
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20076 34354 20132 34366
rect 20076 34302 20078 34354
rect 20130 34302 20132 34354
rect 19852 34242 19908 34254
rect 19852 34190 19854 34242
rect 19906 34190 19908 34242
rect 19628 34076 19796 34132
rect 19516 34020 19572 34030
rect 19516 33926 19572 33964
rect 19628 33906 19684 33918
rect 19628 33854 19630 33906
rect 19682 33854 19684 33906
rect 19516 33460 19572 33470
rect 19516 33122 19572 33404
rect 19516 33070 19518 33122
rect 19570 33070 19572 33122
rect 19516 32228 19572 33070
rect 19628 32340 19684 33854
rect 19740 33236 19796 34076
rect 19852 33460 19908 34190
rect 20076 33684 20132 34302
rect 20412 34132 20468 34524
rect 20076 33618 20132 33628
rect 20300 34130 20468 34132
rect 20300 34078 20414 34130
rect 20466 34078 20468 34130
rect 20300 34076 20468 34078
rect 19852 33394 19908 33404
rect 20300 33458 20356 34076
rect 20412 34066 20468 34076
rect 20300 33406 20302 33458
rect 20354 33406 20356 33458
rect 20300 33394 20356 33406
rect 19740 33180 20132 33236
rect 20076 33124 20132 33180
rect 20076 33068 20244 33124
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32788 20244 33068
rect 19628 32274 19684 32284
rect 20076 32732 20244 32788
rect 19516 32162 19572 32172
rect 19964 32004 20020 32014
rect 19852 31780 19908 31790
rect 19516 31778 19908 31780
rect 19516 31726 19854 31778
rect 19906 31726 19908 31778
rect 19516 31724 19908 31726
rect 19516 30772 19572 31724
rect 19852 31714 19908 31724
rect 19628 31554 19684 31566
rect 19628 31502 19630 31554
rect 19682 31502 19684 31554
rect 19628 31332 19684 31502
rect 19740 31556 19796 31566
rect 19964 31556 20020 31948
rect 20076 31668 20132 32732
rect 20412 32116 20468 32126
rect 20524 32116 20580 35758
rect 20636 35700 20692 36206
rect 20636 35634 20692 35644
rect 20748 36036 20804 36046
rect 20748 35476 20804 35980
rect 20860 35924 20916 36428
rect 20860 35830 20916 35868
rect 21308 36260 21364 36270
rect 20972 35700 21028 35710
rect 20972 35606 21028 35644
rect 20748 34914 20804 35420
rect 21308 35252 21364 36204
rect 20748 34862 20750 34914
rect 20802 34862 20804 34914
rect 20748 34850 20804 34862
rect 20972 34916 21028 34926
rect 20972 34130 21028 34860
rect 20972 34078 20974 34130
rect 21026 34078 21028 34130
rect 20972 34020 21028 34078
rect 21196 34132 21252 34142
rect 21196 34038 21252 34076
rect 20972 33954 21028 33964
rect 20748 33908 20804 33918
rect 20748 33458 20804 33852
rect 20972 33684 21028 33694
rect 20748 33406 20750 33458
rect 20802 33406 20804 33458
rect 20748 33394 20804 33406
rect 20860 33628 20972 33684
rect 20468 32060 20580 32116
rect 20636 32900 20692 32910
rect 20412 31890 20468 32060
rect 20412 31838 20414 31890
rect 20466 31838 20468 31890
rect 20188 31780 20244 31790
rect 20188 31686 20244 31724
rect 20076 31602 20132 31612
rect 19740 31554 20020 31556
rect 19740 31502 19742 31554
rect 19794 31502 20020 31554
rect 19740 31500 20020 31502
rect 20300 31556 20356 31566
rect 19740 31490 19796 31500
rect 20300 31462 20356 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19628 31266 19684 31276
rect 20076 31108 20132 31118
rect 20076 31014 20132 31052
rect 20300 31108 20356 31118
rect 20412 31108 20468 31838
rect 20300 31106 20468 31108
rect 20300 31054 20302 31106
rect 20354 31054 20468 31106
rect 20300 31052 20468 31054
rect 20300 31042 20356 31052
rect 20636 30994 20692 32844
rect 20748 31778 20804 31790
rect 20748 31726 20750 31778
rect 20802 31726 20804 31778
rect 20748 31668 20804 31726
rect 20748 31602 20804 31612
rect 20636 30942 20638 30994
rect 20690 30942 20692 30994
rect 20636 30930 20692 30942
rect 20860 30996 20916 33628
rect 20972 33618 21028 33628
rect 21308 32116 21364 35196
rect 21420 34132 21476 37436
rect 21532 37266 21588 37278
rect 21532 37214 21534 37266
rect 21586 37214 21588 37266
rect 21532 36932 21588 37214
rect 21868 37156 21924 37774
rect 21756 37100 21924 37156
rect 22092 37604 22148 37614
rect 21644 36932 21700 36942
rect 21532 36876 21644 36932
rect 21644 36866 21700 36876
rect 21532 36258 21588 36270
rect 21532 36206 21534 36258
rect 21586 36206 21588 36258
rect 21532 36036 21588 36206
rect 21532 34804 21588 35980
rect 21756 35364 21812 37100
rect 22092 37044 22148 37548
rect 21756 35298 21812 35308
rect 21868 36988 22148 37044
rect 21644 34804 21700 34814
rect 21532 34802 21700 34804
rect 21532 34750 21646 34802
rect 21698 34750 21700 34802
rect 21532 34748 21700 34750
rect 21420 32676 21476 34076
rect 21644 34020 21700 34748
rect 21532 33348 21588 33358
rect 21532 33254 21588 33292
rect 21644 33012 21700 33964
rect 21868 34242 21924 36988
rect 21980 36260 22036 36270
rect 21980 36166 22036 36204
rect 21868 34190 21870 34242
rect 21922 34190 21924 34242
rect 21644 32946 21700 32956
rect 21756 33908 21812 33918
rect 21420 32620 21588 32676
rect 21308 32050 21364 32060
rect 21420 32450 21476 32462
rect 21420 32398 21422 32450
rect 21474 32398 21476 32450
rect 21420 32004 21476 32398
rect 21420 31938 21476 31948
rect 21420 31554 21476 31566
rect 21420 31502 21422 31554
rect 21474 31502 21476 31554
rect 21420 31444 21476 31502
rect 21420 31378 21476 31388
rect 21532 31332 21588 32620
rect 21644 32562 21700 32574
rect 21644 32510 21646 32562
rect 21698 32510 21700 32562
rect 21644 32004 21700 32510
rect 21644 31938 21700 31948
rect 21532 31276 21700 31332
rect 20972 31220 21028 31230
rect 20972 31218 21588 31220
rect 20972 31166 20974 31218
rect 21026 31166 21588 31218
rect 20972 31164 21588 31166
rect 20972 31154 21028 31164
rect 20860 30940 21028 30996
rect 19516 30706 19572 30716
rect 19628 30882 19684 30894
rect 19628 30830 19630 30882
rect 19682 30830 19684 30882
rect 19628 30324 19684 30830
rect 19404 30268 19572 30324
rect 19292 30158 19294 30210
rect 19346 30158 19348 30210
rect 19292 29988 19348 30158
rect 19292 29922 19348 29932
rect 19404 30100 19460 30110
rect 19404 29652 19460 30044
rect 19516 29988 19572 30268
rect 19628 30258 19684 30268
rect 19964 30772 20020 30782
rect 19964 30436 20020 30716
rect 19964 30210 20020 30380
rect 19964 30158 19966 30210
rect 20018 30158 20020 30210
rect 19964 30100 20020 30158
rect 20860 30770 20916 30782
rect 20860 30718 20862 30770
rect 20914 30718 20916 30770
rect 20860 30660 20916 30718
rect 19964 30034 20020 30044
rect 20412 30100 20468 30110
rect 20412 30006 20468 30044
rect 19516 29932 19684 29988
rect 19516 29652 19572 29662
rect 19404 29596 19516 29652
rect 19516 29558 19572 29596
rect 19292 29092 19348 29102
rect 19292 28644 19348 29036
rect 19292 28550 19348 28588
rect 19628 27972 19684 29932
rect 20860 29876 20916 30604
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20860 29810 20916 29820
rect 19836 29754 20100 29764
rect 19740 29652 19796 29662
rect 19740 29426 19796 29596
rect 20076 29652 20132 29662
rect 20860 29652 20916 29662
rect 20972 29652 21028 30940
rect 21420 30882 21476 30894
rect 21420 30830 21422 30882
rect 21474 30830 21476 30882
rect 21420 30772 21476 30830
rect 21420 30706 21476 30716
rect 21196 30212 21252 30222
rect 20076 29558 20132 29596
rect 20412 29650 21140 29652
rect 20412 29598 20862 29650
rect 20914 29598 21140 29650
rect 20412 29596 21140 29598
rect 20412 29538 20468 29596
rect 20860 29586 20916 29596
rect 20412 29486 20414 29538
rect 20466 29486 20468 29538
rect 20412 29474 20468 29486
rect 19740 29374 19742 29426
rect 19794 29374 19796 29426
rect 19740 29362 19796 29374
rect 19964 29426 20020 29438
rect 19964 29374 19966 29426
rect 20018 29374 20020 29426
rect 19964 29316 20020 29374
rect 20188 29428 20244 29438
rect 20244 29372 20356 29428
rect 20188 29334 20244 29372
rect 19964 29250 20020 29260
rect 20076 28756 20132 28766
rect 20132 28700 20244 28756
rect 20076 28662 20132 28700
rect 20188 28532 20244 28700
rect 20300 28644 20356 29372
rect 20748 29316 20804 29326
rect 20412 28644 20468 28654
rect 20300 28642 20468 28644
rect 20300 28590 20414 28642
rect 20466 28590 20468 28642
rect 20300 28588 20468 28590
rect 20412 28578 20468 28588
rect 20748 28642 20804 29260
rect 20748 28590 20750 28642
rect 20802 28590 20804 28642
rect 20748 28578 20804 28590
rect 20188 28476 20356 28532
rect 20300 28420 20356 28476
rect 20524 28420 20580 28430
rect 20300 28418 20580 28420
rect 20300 28366 20526 28418
rect 20578 28366 20580 28418
rect 20300 28364 20580 28366
rect 20524 28354 20580 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 28196 20244 28206
rect 19628 27878 19684 27916
rect 19404 27858 19460 27870
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 19404 27524 19460 27806
rect 19404 27186 19460 27468
rect 19404 27134 19406 27186
rect 19458 27134 19460 27186
rect 19404 27122 19460 27134
rect 19964 27858 20020 27870
rect 19964 27806 19966 27858
rect 20018 27806 20020 27858
rect 19964 27076 20020 27806
rect 20188 27186 20244 28140
rect 20636 27972 20692 27982
rect 20636 27878 20692 27916
rect 20972 27970 21028 27982
rect 20972 27918 20974 27970
rect 21026 27918 21028 27970
rect 20188 27134 20190 27186
rect 20242 27134 20244 27186
rect 20188 27122 20244 27134
rect 19964 27010 20020 27020
rect 20972 26908 21028 27918
rect 18956 26852 19124 26908
rect 19292 26852 19348 26862
rect 17948 26460 18228 26516
rect 17836 26238 17838 26290
rect 17890 26238 17892 26290
rect 17836 26068 17892 26238
rect 17388 25454 17390 25506
rect 17442 25454 17444 25506
rect 17388 25442 17444 25454
rect 17500 26012 17892 26068
rect 17948 26292 18004 26302
rect 17388 25060 17444 25070
rect 17500 25060 17556 26012
rect 17724 25620 17780 25630
rect 17948 25620 18004 26236
rect 17724 25618 18004 25620
rect 17724 25566 17726 25618
rect 17778 25566 18004 25618
rect 17724 25564 18004 25566
rect 17612 25394 17668 25406
rect 17612 25342 17614 25394
rect 17666 25342 17668 25394
rect 17612 25172 17668 25342
rect 17724 25284 17780 25564
rect 18172 25508 18228 26460
rect 18956 26404 19012 26852
rect 18956 26348 19236 26404
rect 18508 26292 18564 26302
rect 18508 26198 18564 26236
rect 19068 26178 19124 26190
rect 19068 26126 19070 26178
rect 19122 26126 19124 26178
rect 17724 25218 17780 25228
rect 17836 25506 18228 25508
rect 17836 25454 18174 25506
rect 18226 25454 18228 25506
rect 17836 25452 18228 25454
rect 17612 25106 17668 25116
rect 17444 25004 17556 25060
rect 17388 24994 17444 25004
rect 17612 24948 17668 24958
rect 17836 24948 17892 25452
rect 18172 25442 18228 25452
rect 18508 25508 18564 25518
rect 17612 24946 17892 24948
rect 17612 24894 17614 24946
rect 17666 24894 17892 24946
rect 17612 24892 17892 24894
rect 17948 25172 18004 25182
rect 17612 24882 17668 24892
rect 17164 24770 17220 24780
rect 17836 24724 17892 24734
rect 17836 24630 17892 24668
rect 16828 24546 16884 24556
rect 17948 23938 18004 25116
rect 17948 23886 17950 23938
rect 18002 23886 18004 23938
rect 17948 23874 18004 23886
rect 16940 23828 16996 23838
rect 16604 23826 16996 23828
rect 16604 23774 16942 23826
rect 16994 23774 16996 23826
rect 16604 23772 16996 23774
rect 16156 23378 16212 23436
rect 16156 23326 16158 23378
rect 16210 23326 16212 23378
rect 16156 23314 16212 23326
rect 16492 23380 16548 23772
rect 16940 23762 16996 23772
rect 18172 23828 18228 23838
rect 18508 23828 18564 25452
rect 18844 25506 18900 25518
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 25396 18900 25454
rect 18844 25330 18900 25340
rect 18620 25284 18676 25294
rect 18620 24276 18676 25228
rect 19068 25284 19124 26126
rect 19068 25218 19124 25228
rect 19180 24610 19236 26348
rect 19292 25506 19348 26796
rect 20412 26852 20468 26862
rect 19836 26684 20100 26694
rect 19516 26628 19572 26638
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19516 26516 19572 26572
rect 19516 26514 19908 26516
rect 19516 26462 19518 26514
rect 19570 26462 19908 26514
rect 19516 26460 19908 26462
rect 19516 26450 19572 26460
rect 19852 25620 19908 26460
rect 20412 26514 20468 26796
rect 20412 26462 20414 26514
rect 20466 26462 20468 26514
rect 19964 26178 20020 26190
rect 19964 26126 19966 26178
rect 20018 26126 20020 26178
rect 19964 26068 20020 26126
rect 19964 26002 20020 26012
rect 20412 25956 20468 26462
rect 20412 25890 20468 25900
rect 20636 26852 21028 26908
rect 21084 26908 21140 29596
rect 21196 29426 21252 30156
rect 21532 30210 21588 31164
rect 21532 30158 21534 30210
rect 21586 30158 21588 30210
rect 21532 30146 21588 30158
rect 21644 30212 21700 31276
rect 21756 30436 21812 33852
rect 21868 32900 21924 34190
rect 22092 35028 22148 35038
rect 21980 33572 22036 33582
rect 21980 33236 22036 33516
rect 21980 33142 22036 33180
rect 21868 32834 21924 32844
rect 21868 32674 21924 32686
rect 21868 32622 21870 32674
rect 21922 32622 21924 32674
rect 21868 31780 21924 32622
rect 21868 31714 21924 31724
rect 21980 32564 22036 32574
rect 21868 30882 21924 30894
rect 21868 30830 21870 30882
rect 21922 30830 21924 30882
rect 21868 30660 21924 30830
rect 21868 30594 21924 30604
rect 21868 30436 21924 30446
rect 21756 30434 21924 30436
rect 21756 30382 21870 30434
rect 21922 30382 21924 30434
rect 21756 30380 21924 30382
rect 21868 30370 21924 30380
rect 21980 30436 22036 32508
rect 21980 30370 22036 30380
rect 21756 30212 21812 30222
rect 21644 30210 21812 30212
rect 21644 30158 21758 30210
rect 21810 30158 21812 30210
rect 21644 30156 21812 30158
rect 22092 30212 22148 34972
rect 22204 34130 22260 34142
rect 22204 34078 22206 34130
rect 22258 34078 22260 34130
rect 22204 33124 22260 34078
rect 22316 33460 22372 43484
rect 22428 41970 22484 45388
rect 22764 45106 22820 45612
rect 22988 45220 23044 48300
rect 23436 48354 23492 48366
rect 23436 48302 23438 48354
rect 23490 48302 23492 48354
rect 23100 48244 23156 48254
rect 23324 48244 23380 48254
rect 23100 48242 23380 48244
rect 23100 48190 23102 48242
rect 23154 48190 23326 48242
rect 23378 48190 23380 48242
rect 23100 48188 23380 48190
rect 23100 48178 23156 48188
rect 23324 48178 23380 48188
rect 23436 48244 23492 48302
rect 23436 48178 23492 48188
rect 23100 46676 23156 46686
rect 23100 46582 23156 46620
rect 23548 46676 23604 51436
rect 23772 50428 23828 53452
rect 23996 52948 24052 53454
rect 24444 53508 24500 53678
rect 24444 53442 24500 53452
rect 24780 53506 24836 54348
rect 25116 53844 25172 53854
rect 25116 53730 25172 53788
rect 25116 53678 25118 53730
rect 25170 53678 25172 53730
rect 25116 53666 25172 53678
rect 24780 53454 24782 53506
rect 24834 53454 24836 53506
rect 24780 53442 24836 53454
rect 24892 53618 24948 53630
rect 24892 53566 24894 53618
rect 24946 53566 24948 53618
rect 24892 53508 24948 53566
rect 23996 52882 24052 52892
rect 24780 52724 24836 52734
rect 24892 52724 24948 53452
rect 24836 52668 24948 52724
rect 25116 52722 25172 52734
rect 25116 52670 25118 52722
rect 25170 52670 25172 52722
rect 24780 52658 24836 52668
rect 25116 50820 25172 52670
rect 25228 52388 25284 54462
rect 25340 53508 25396 55022
rect 27580 55076 27636 55086
rect 27580 54982 27636 55020
rect 26012 54404 26068 54414
rect 26012 54310 26068 54348
rect 28140 54402 28196 54414
rect 28140 54350 28142 54402
rect 28194 54350 28196 54402
rect 26348 53844 26404 53854
rect 26348 53750 26404 53788
rect 26572 53844 26628 53854
rect 25564 53508 25620 53518
rect 25340 53452 25564 53508
rect 25564 53414 25620 53452
rect 26236 53506 26292 53518
rect 26236 53454 26238 53506
rect 26290 53454 26292 53506
rect 25452 52948 25508 52958
rect 25340 52892 25452 52948
rect 25340 52722 25396 52892
rect 25452 52854 25508 52892
rect 25900 52946 25956 52958
rect 25900 52894 25902 52946
rect 25954 52894 25956 52946
rect 25340 52670 25342 52722
rect 25394 52670 25396 52722
rect 25340 52658 25396 52670
rect 25228 52164 25284 52332
rect 25228 51380 25284 52108
rect 25452 52052 25508 52062
rect 25340 51380 25396 51390
rect 25228 51378 25396 51380
rect 25228 51326 25342 51378
rect 25394 51326 25396 51378
rect 25228 51324 25396 51326
rect 25340 51314 25396 51324
rect 25116 50764 25284 50820
rect 24220 50706 24276 50718
rect 24220 50654 24222 50706
rect 24274 50654 24276 50706
rect 23772 50372 24164 50428
rect 24108 49700 24164 50372
rect 24220 50148 24276 50654
rect 24892 50652 25172 50708
rect 24556 50596 24612 50606
rect 24556 50370 24612 50540
rect 24780 50484 24836 50494
rect 24892 50484 24948 50652
rect 24780 50482 24948 50484
rect 24780 50430 24782 50482
rect 24834 50430 24948 50482
rect 24780 50428 24948 50430
rect 25116 50428 25172 50652
rect 25228 50594 25284 50764
rect 25228 50542 25230 50594
rect 25282 50542 25284 50594
rect 25228 50530 25284 50542
rect 25452 50596 25508 51996
rect 25900 51268 25956 52894
rect 26124 52948 26180 52958
rect 26236 52948 26292 53454
rect 26460 53508 26516 53518
rect 26572 53508 26628 53788
rect 28140 53844 28196 54350
rect 28140 53778 28196 53788
rect 26460 53506 26628 53508
rect 26460 53454 26462 53506
rect 26514 53454 26628 53506
rect 26460 53452 26628 53454
rect 26460 53442 26516 53452
rect 26124 52946 26292 52948
rect 26124 52894 26126 52946
rect 26178 52894 26292 52946
rect 26124 52892 26292 52894
rect 26124 52882 26180 52892
rect 25900 51202 25956 51212
rect 26012 52834 26068 52846
rect 26012 52782 26014 52834
rect 26066 52782 26068 52834
rect 25452 50482 25508 50540
rect 26012 50596 26068 52782
rect 26236 52052 26292 52892
rect 26236 51986 26292 51996
rect 26460 52612 26516 52622
rect 26460 52052 26516 52556
rect 26460 51986 26516 51996
rect 26124 51268 26180 51278
rect 26124 51266 26516 51268
rect 26124 51214 26126 51266
rect 26178 51214 26516 51266
rect 26124 51212 26516 51214
rect 26124 51202 26180 51212
rect 26460 50706 26516 51212
rect 26460 50654 26462 50706
rect 26514 50654 26516 50706
rect 26460 50642 26516 50654
rect 26012 50530 26068 50540
rect 26236 50594 26292 50606
rect 26236 50542 26238 50594
rect 26290 50542 26292 50594
rect 25452 50430 25454 50482
rect 25506 50430 25508 50482
rect 24556 50318 24558 50370
rect 24610 50318 24612 50370
rect 24556 50306 24612 50318
rect 24668 50372 24724 50382
rect 24668 50278 24724 50316
rect 24780 50148 24836 50428
rect 25116 50372 25284 50428
rect 25452 50418 25508 50430
rect 24220 50092 24836 50148
rect 25228 49922 25284 50372
rect 25228 49870 25230 49922
rect 25282 49870 25284 49922
rect 25228 49858 25284 49870
rect 25788 50370 25844 50382
rect 25788 50318 25790 50370
rect 25842 50318 25844 50370
rect 25788 49700 25844 50318
rect 26236 50260 26292 50542
rect 26572 50428 26628 53452
rect 26684 53506 26740 53518
rect 26684 53454 26686 53506
rect 26738 53454 26740 53506
rect 26684 53058 26740 53454
rect 26684 53006 26686 53058
rect 26738 53006 26740 53058
rect 26684 52948 26740 53006
rect 26684 52882 26740 52892
rect 27020 52948 27076 52958
rect 27020 52836 27076 52892
rect 27468 52836 27524 52846
rect 27020 52834 27636 52836
rect 27020 52782 27470 52834
rect 27522 52782 27636 52834
rect 27020 52780 27636 52782
rect 27468 52770 27524 52780
rect 27020 52276 27076 52286
rect 27020 52164 27076 52220
rect 27468 52164 27524 52174
rect 27020 52162 27524 52164
rect 27020 52110 27022 52162
rect 27074 52110 27470 52162
rect 27522 52110 27524 52162
rect 27020 52108 27524 52110
rect 27020 52098 27076 52108
rect 26684 52052 26740 52062
rect 26684 50708 26740 51996
rect 26684 50594 26740 50652
rect 27356 50708 27412 50718
rect 27356 50614 27412 50652
rect 26684 50542 26686 50594
rect 26738 50542 26740 50594
rect 26684 50530 26740 50542
rect 26796 50596 26852 50606
rect 26796 50502 26852 50540
rect 26236 50194 26292 50204
rect 26460 50372 26628 50428
rect 24108 49644 24612 49700
rect 24332 49476 24388 49486
rect 23884 48468 23940 48478
rect 23884 48354 23940 48412
rect 23884 48302 23886 48354
rect 23938 48302 23940 48354
rect 23884 48290 23940 48302
rect 23996 48354 24052 48366
rect 23996 48302 23998 48354
rect 24050 48302 24052 48354
rect 23660 48244 23716 48254
rect 23996 48244 24052 48302
rect 23660 48242 23828 48244
rect 23660 48190 23662 48242
rect 23714 48190 23828 48242
rect 23660 48188 23828 48190
rect 23660 48178 23716 48188
rect 23548 46610 23604 46620
rect 23660 46562 23716 46574
rect 23660 46510 23662 46562
rect 23714 46510 23716 46562
rect 23660 46452 23716 46510
rect 23660 46386 23716 46396
rect 23660 45778 23716 45790
rect 23660 45726 23662 45778
rect 23714 45726 23716 45778
rect 23324 45332 23380 45342
rect 23324 45238 23380 45276
rect 22988 45154 23044 45164
rect 22764 45054 22766 45106
rect 22818 45054 22820 45106
rect 22764 45042 22820 45054
rect 23660 44996 23716 45726
rect 23660 44930 23716 44940
rect 22988 44884 23044 44894
rect 22764 44882 23044 44884
rect 22764 44830 22990 44882
rect 23042 44830 23044 44882
rect 22764 44828 23044 44830
rect 22652 44436 22708 44446
rect 22652 44098 22708 44380
rect 22652 44046 22654 44098
rect 22706 44046 22708 44098
rect 22652 42868 22708 44046
rect 22652 42802 22708 42812
rect 22428 41918 22430 41970
rect 22482 41918 22484 41970
rect 22428 41906 22484 41918
rect 22540 42756 22596 42766
rect 22428 39506 22484 39518
rect 22428 39454 22430 39506
rect 22482 39454 22484 39506
rect 22428 38836 22484 39454
rect 22428 38770 22484 38780
rect 22540 38668 22596 42700
rect 22652 40628 22708 40638
rect 22652 40534 22708 40572
rect 22764 40068 22820 44828
rect 22988 44818 23044 44828
rect 23100 44772 23156 44782
rect 23100 44324 23156 44716
rect 22988 44322 23156 44324
rect 22988 44270 23102 44322
rect 23154 44270 23156 44322
rect 22988 44268 23156 44270
rect 22876 43540 22932 43550
rect 22876 42756 22932 43484
rect 22876 42690 22932 42700
rect 22876 41860 22932 41870
rect 22876 41766 22932 41804
rect 22876 41300 22932 41310
rect 22876 41206 22932 41244
rect 22428 38612 22596 38668
rect 22652 40012 22820 40068
rect 22428 37940 22484 38612
rect 22428 37846 22484 37884
rect 22540 37380 22596 37390
rect 22540 36482 22596 37324
rect 22652 37156 22708 40012
rect 22988 39956 23044 44268
rect 23100 44258 23156 44268
rect 23436 44434 23492 44446
rect 23436 44382 23438 44434
rect 23490 44382 23492 44434
rect 23436 43988 23492 44382
rect 23436 43922 23492 43932
rect 23436 43538 23492 43550
rect 23436 43486 23438 43538
rect 23490 43486 23492 43538
rect 23100 43426 23156 43438
rect 23100 43374 23102 43426
rect 23154 43374 23156 43426
rect 23100 43204 23156 43374
rect 23100 43138 23156 43148
rect 23100 42532 23156 42542
rect 23436 42532 23492 43486
rect 23100 42530 23492 42532
rect 23100 42478 23102 42530
rect 23154 42478 23492 42530
rect 23100 42476 23492 42478
rect 23100 42084 23156 42476
rect 23772 42308 23828 48188
rect 23996 48178 24052 48188
rect 23884 48132 23940 48142
rect 23884 42756 23940 48076
rect 23996 48018 24052 48030
rect 23996 47966 23998 48018
rect 24050 47966 24052 48018
rect 23996 46340 24052 47966
rect 24220 46676 24276 46686
rect 24220 46582 24276 46620
rect 24108 46340 24164 46350
rect 23996 46284 24108 46340
rect 24108 46274 24164 46284
rect 24332 46228 24388 49420
rect 24556 49138 24612 49644
rect 25788 49606 25844 49644
rect 24556 49086 24558 49138
rect 24610 49086 24612 49138
rect 24556 49074 24612 49086
rect 25340 49586 25396 49598
rect 25340 49534 25342 49586
rect 25394 49534 25396 49586
rect 24668 49028 24724 49038
rect 24668 48934 24724 48972
rect 25340 48580 25396 49534
rect 25676 49026 25732 49038
rect 25676 48974 25678 49026
rect 25730 48974 25732 49026
rect 25340 48514 25396 48524
rect 25452 48914 25508 48926
rect 25452 48862 25454 48914
rect 25506 48862 25508 48914
rect 24556 48244 24612 48254
rect 24556 48150 24612 48188
rect 25452 47572 25508 48862
rect 25452 47506 25508 47516
rect 25564 47458 25620 47470
rect 25564 47406 25566 47458
rect 25618 47406 25620 47458
rect 25564 47348 25620 47406
rect 25564 47282 25620 47292
rect 25228 46676 25284 46686
rect 25228 46582 25284 46620
rect 24220 46172 24388 46228
rect 24780 46562 24836 46574
rect 24780 46510 24782 46562
rect 24834 46510 24836 46562
rect 24220 46004 24276 46172
rect 24780 46116 24836 46510
rect 24108 45948 24276 46004
rect 24332 46060 24836 46116
rect 24892 46340 24948 46350
rect 23996 44660 24052 44670
rect 23996 43538 24052 44604
rect 23996 43486 23998 43538
rect 24050 43486 24052 43538
rect 23996 43474 24052 43486
rect 23884 42690 23940 42700
rect 23884 42532 23940 42542
rect 23884 42530 24052 42532
rect 23884 42478 23886 42530
rect 23938 42478 24052 42530
rect 23884 42476 24052 42478
rect 23884 42466 23940 42476
rect 23772 42252 23940 42308
rect 23100 42018 23156 42028
rect 23436 41972 23492 41982
rect 23212 41860 23268 41870
rect 23100 41858 23268 41860
rect 23100 41806 23214 41858
rect 23266 41806 23268 41858
rect 23100 41804 23268 41806
rect 23100 41748 23156 41804
rect 23212 41794 23268 41804
rect 23100 40740 23156 41692
rect 23100 40674 23156 40684
rect 23212 41188 23268 41198
rect 23212 40628 23268 41132
rect 23212 40562 23268 40572
rect 23436 40628 23492 41916
rect 23436 40562 23492 40572
rect 23772 41074 23828 41086
rect 23772 41022 23774 41074
rect 23826 41022 23828 41074
rect 23100 40404 23156 40414
rect 23100 40310 23156 40348
rect 23772 40404 23828 41022
rect 23772 40338 23828 40348
rect 22876 39900 23044 39956
rect 23772 40178 23828 40190
rect 23772 40126 23774 40178
rect 23826 40126 23828 40178
rect 22764 38722 22820 38734
rect 22764 38670 22766 38722
rect 22818 38670 22820 38722
rect 22764 37604 22820 38670
rect 22764 37538 22820 37548
rect 22876 38724 22932 39900
rect 22988 39732 23044 39742
rect 22988 39730 23380 39732
rect 22988 39678 22990 39730
rect 23042 39678 23380 39730
rect 22988 39676 23380 39678
rect 22988 39172 23044 39676
rect 23324 39618 23380 39676
rect 23324 39566 23326 39618
rect 23378 39566 23380 39618
rect 23324 39554 23380 39566
rect 22988 39106 23044 39116
rect 23772 39058 23828 40126
rect 23884 39506 23940 42252
rect 23996 41972 24052 42476
rect 23996 41188 24052 41916
rect 23996 41122 24052 41132
rect 24108 40626 24164 45948
rect 24220 45780 24276 45790
rect 24332 45780 24388 46060
rect 24220 45778 24388 45780
rect 24220 45726 24222 45778
rect 24274 45726 24388 45778
rect 24220 45724 24388 45726
rect 24220 45714 24276 45724
rect 24332 44098 24388 45724
rect 24444 45890 24500 45902
rect 24444 45838 24446 45890
rect 24498 45838 24500 45890
rect 24444 44660 24500 45838
rect 24780 45890 24836 45902
rect 24780 45838 24782 45890
rect 24834 45838 24836 45890
rect 24556 45780 24612 45790
rect 24556 45686 24612 45724
rect 24668 44996 24724 45006
rect 24668 44902 24724 44940
rect 24444 44594 24500 44604
rect 24668 44436 24724 44446
rect 24780 44436 24836 45838
rect 24892 45778 24948 46284
rect 24892 45726 24894 45778
rect 24946 45726 24948 45778
rect 24892 45714 24948 45726
rect 25340 44996 25396 45006
rect 25340 44902 25396 44940
rect 25116 44660 25172 44670
rect 25172 44604 25284 44660
rect 25116 44594 25172 44604
rect 24780 44380 25060 44436
rect 24668 44212 24724 44380
rect 24780 44212 24836 44222
rect 24668 44156 24780 44212
rect 24780 44118 24836 44156
rect 24332 44046 24334 44098
rect 24386 44046 24388 44098
rect 24332 43988 24388 44046
rect 24332 43092 24388 43932
rect 24668 43540 24724 43550
rect 24668 43446 24724 43484
rect 24332 43026 24388 43036
rect 24668 42980 24724 42990
rect 24668 42886 24724 42924
rect 24556 42642 24612 42654
rect 24556 42590 24558 42642
rect 24610 42590 24612 42642
rect 24332 42530 24388 42542
rect 24332 42478 24334 42530
rect 24386 42478 24388 42530
rect 24332 41300 24388 42478
rect 24556 41972 24612 42590
rect 24556 41906 24612 41916
rect 24668 42530 24724 42542
rect 24668 42478 24670 42530
rect 24722 42478 24724 42530
rect 24668 41300 24724 42478
rect 24780 41972 24836 41982
rect 24780 41878 24836 41916
rect 24780 41300 24836 41310
rect 24668 41244 24780 41300
rect 24836 41244 24948 41300
rect 24332 41234 24388 41244
rect 24780 41234 24836 41244
rect 24892 41186 24948 41244
rect 25004 41298 25060 44380
rect 25228 44324 25284 44604
rect 25228 44230 25284 44268
rect 25116 44212 25172 44222
rect 25116 44118 25172 44156
rect 25676 43708 25732 48974
rect 26460 48354 26516 50372
rect 27468 49476 27524 52108
rect 27580 51940 27636 52780
rect 27580 51884 28084 51940
rect 27580 51268 27636 51278
rect 27580 49922 27636 51212
rect 27580 49870 27582 49922
rect 27634 49870 27636 49922
rect 27580 49858 27636 49870
rect 27692 49586 27748 49598
rect 27692 49534 27694 49586
rect 27746 49534 27748 49586
rect 27468 49420 27636 49476
rect 27132 49028 27188 49038
rect 27132 48934 27188 48972
rect 27356 48914 27412 48926
rect 27356 48862 27358 48914
rect 27410 48862 27412 48914
rect 27356 48692 27412 48862
rect 27356 48626 27412 48636
rect 27468 48580 27524 48590
rect 26460 48302 26462 48354
rect 26514 48302 26516 48354
rect 26460 48290 26516 48302
rect 27356 48354 27412 48366
rect 27356 48302 27358 48354
rect 27410 48302 27412 48354
rect 26572 48244 26628 48254
rect 26572 48150 26628 48188
rect 27132 48242 27188 48254
rect 27132 48190 27134 48242
rect 27186 48190 27188 48242
rect 26908 47572 26964 47582
rect 25788 47348 25844 47358
rect 25788 47346 26068 47348
rect 25788 47294 25790 47346
rect 25842 47294 26068 47346
rect 25788 47292 26068 47294
rect 25788 47282 25844 47292
rect 25900 45220 25956 45230
rect 25788 44996 25844 45006
rect 25788 44902 25844 44940
rect 25788 44660 25844 44670
rect 25788 44434 25844 44604
rect 25788 44382 25790 44434
rect 25842 44382 25844 44434
rect 25788 44370 25844 44382
rect 25676 43652 25844 43708
rect 25564 43538 25620 43550
rect 25564 43486 25566 43538
rect 25618 43486 25620 43538
rect 25004 41246 25006 41298
rect 25058 41246 25060 41298
rect 25004 41234 25060 41246
rect 25116 43428 25172 43438
rect 25340 43428 25396 43438
rect 24892 41134 24894 41186
rect 24946 41134 24948 41186
rect 24892 41122 24948 41134
rect 24108 40574 24110 40626
rect 24162 40574 24164 40626
rect 24108 40178 24164 40574
rect 24780 41076 24836 41086
rect 24780 40516 24836 41020
rect 24780 40450 24836 40460
rect 24108 40126 24110 40178
rect 24162 40126 24164 40178
rect 24108 40114 24164 40126
rect 25004 40180 25060 40190
rect 23884 39454 23886 39506
rect 23938 39454 23940 39506
rect 23884 39442 23940 39454
rect 24668 39844 24724 39854
rect 23772 39006 23774 39058
rect 23826 39006 23828 39058
rect 23324 38836 23380 38846
rect 23212 38724 23268 38734
rect 22876 38722 23268 38724
rect 22876 38670 23214 38722
rect 23266 38670 23268 38722
rect 22876 38668 23268 38670
rect 22764 37268 22820 37278
rect 22876 37268 22932 38668
rect 23212 38658 23268 38668
rect 23212 38052 23268 38062
rect 22988 37826 23044 37838
rect 22988 37774 22990 37826
rect 23042 37774 23044 37826
rect 22988 37380 23044 37774
rect 22988 37314 23044 37324
rect 23100 37604 23156 37614
rect 22764 37266 22932 37268
rect 22764 37214 22766 37266
rect 22818 37214 22932 37266
rect 22764 37212 22932 37214
rect 22764 37202 22820 37212
rect 22652 37090 22708 37100
rect 23100 37156 23156 37548
rect 23100 37090 23156 37100
rect 22540 36430 22542 36482
rect 22594 36430 22596 36482
rect 22540 36418 22596 36430
rect 22876 36372 22932 36382
rect 22876 36278 22932 36316
rect 22876 35924 22932 35934
rect 22876 35810 22932 35868
rect 22876 35758 22878 35810
rect 22930 35758 22932 35810
rect 22876 35746 22932 35758
rect 22540 35700 22596 35710
rect 22540 34914 22596 35644
rect 22540 34862 22542 34914
rect 22594 34862 22596 34914
rect 22540 33460 22596 34862
rect 22988 35698 23044 35710
rect 22988 35646 22990 35698
rect 23042 35646 23044 35698
rect 22764 34804 22820 34814
rect 22652 34692 22708 34702
rect 22652 34130 22708 34636
rect 22764 34692 22820 34748
rect 22988 34692 23044 35646
rect 23212 35586 23268 37996
rect 23212 35534 23214 35586
rect 23266 35534 23268 35586
rect 23212 35522 23268 35534
rect 23324 36932 23380 38780
rect 23772 38668 23828 39006
rect 24668 39058 24724 39788
rect 24668 39006 24670 39058
rect 24722 39006 24724 39058
rect 24220 38948 24276 38958
rect 24220 38854 24276 38892
rect 23772 38612 23940 38668
rect 22764 34690 23044 34692
rect 22764 34638 22766 34690
rect 22818 34638 23044 34690
rect 22764 34636 23044 34638
rect 22764 34626 22820 34636
rect 23324 34580 23380 36876
rect 23436 37826 23492 37838
rect 23436 37774 23438 37826
rect 23490 37774 23492 37826
rect 23436 37716 23492 37774
rect 23436 35476 23492 37660
rect 23772 37826 23828 37838
rect 23772 37774 23774 37826
rect 23826 37774 23828 37826
rect 23660 37268 23716 37278
rect 23436 35410 23492 35420
rect 23548 35698 23604 35710
rect 23548 35646 23550 35698
rect 23602 35646 23604 35698
rect 23548 35028 23604 35646
rect 23660 35252 23716 37212
rect 23660 35186 23716 35196
rect 23772 35140 23828 37774
rect 23884 37716 23940 38612
rect 24108 38050 24164 38062
rect 24108 37998 24110 38050
rect 24162 37998 24164 38050
rect 24108 37828 24164 37998
rect 24668 37940 24724 39006
rect 25004 38052 25060 40124
rect 25116 39058 25172 43372
rect 25228 43426 25396 43428
rect 25228 43374 25342 43426
rect 25394 43374 25396 43426
rect 25228 43372 25396 43374
rect 25228 41972 25284 43372
rect 25340 43362 25396 43372
rect 25452 42866 25508 42878
rect 25452 42814 25454 42866
rect 25506 42814 25508 42866
rect 25452 42308 25508 42814
rect 25452 42242 25508 42252
rect 25228 41916 25396 41972
rect 25340 41858 25396 41916
rect 25340 41806 25342 41858
rect 25394 41806 25396 41858
rect 25340 41794 25396 41806
rect 25564 40628 25620 43486
rect 25676 43538 25732 43550
rect 25676 43486 25678 43538
rect 25730 43486 25732 43538
rect 25676 43204 25732 43486
rect 25676 43138 25732 43148
rect 25676 42754 25732 42766
rect 25676 42702 25678 42754
rect 25730 42702 25732 42754
rect 25676 41972 25732 42702
rect 25676 41878 25732 41916
rect 25788 41636 25844 43652
rect 25900 43538 25956 45164
rect 26012 44546 26068 47292
rect 26908 46002 26964 47516
rect 26908 45950 26910 46002
rect 26962 45950 26964 46002
rect 26908 45938 26964 45950
rect 26796 45890 26852 45902
rect 26796 45838 26798 45890
rect 26850 45838 26852 45890
rect 26236 45218 26292 45230
rect 26236 45166 26238 45218
rect 26290 45166 26292 45218
rect 26124 45108 26180 45118
rect 26124 45014 26180 45052
rect 26236 44548 26292 45166
rect 26012 44494 26014 44546
rect 26066 44494 26068 44546
rect 26012 44482 26068 44494
rect 26124 44492 26292 44548
rect 26348 45220 26404 45230
rect 25900 43486 25902 43538
rect 25954 43486 25956 43538
rect 25900 43474 25956 43486
rect 26124 43428 26180 44492
rect 26236 44324 26292 44334
rect 26236 43428 26292 44268
rect 26348 43650 26404 45164
rect 26796 44436 26852 45838
rect 26348 43598 26350 43650
rect 26402 43598 26404 43650
rect 26348 43586 26404 43598
rect 26460 44380 26852 44436
rect 26348 43428 26404 43438
rect 26236 43372 26348 43428
rect 26124 43362 26180 43372
rect 26348 43362 26404 43372
rect 26236 42642 26292 42654
rect 26236 42590 26238 42642
rect 26290 42590 26292 42642
rect 26236 42420 26292 42590
rect 26236 42354 26292 42364
rect 26348 42308 26404 42318
rect 25788 41570 25844 41580
rect 25900 42084 25956 42094
rect 25900 41858 25956 42028
rect 26348 42084 26404 42252
rect 26348 41990 26404 42028
rect 25900 41806 25902 41858
rect 25954 41806 25956 41858
rect 25900 41076 25956 41806
rect 26236 41972 26292 41982
rect 26236 41412 26292 41916
rect 26236 41346 26292 41356
rect 25900 41010 25956 41020
rect 25676 40628 25732 40638
rect 25564 40626 25732 40628
rect 25564 40574 25678 40626
rect 25730 40574 25732 40626
rect 25564 40572 25732 40574
rect 25676 40562 25732 40572
rect 26124 40404 26180 40414
rect 25452 40402 26180 40404
rect 25452 40350 26126 40402
rect 26178 40350 26180 40402
rect 25452 40348 26180 40350
rect 25340 40180 25396 40190
rect 25340 40086 25396 40124
rect 25452 40068 25508 40348
rect 26124 40338 26180 40348
rect 25452 39844 25508 40012
rect 25452 39778 25508 39788
rect 25564 40178 25620 40190
rect 25564 40126 25566 40178
rect 25618 40126 25620 40178
rect 25564 39508 25620 40126
rect 25564 39442 25620 39452
rect 25676 40180 25732 40190
rect 26348 40180 26404 40190
rect 25676 40178 26404 40180
rect 25676 40126 25678 40178
rect 25730 40126 26350 40178
rect 26402 40126 26404 40178
rect 25676 40124 26404 40126
rect 25116 39006 25118 39058
rect 25170 39006 25172 39058
rect 25116 38994 25172 39006
rect 25564 38724 25620 38762
rect 25564 38658 25620 38668
rect 25004 37996 25284 38052
rect 24108 37762 24164 37772
rect 24444 37884 24724 37940
rect 25228 37940 25284 37996
rect 25228 37938 25396 37940
rect 25228 37886 25230 37938
rect 25282 37886 25396 37938
rect 25228 37884 25396 37886
rect 23884 37650 23940 37660
rect 24444 37492 24500 37884
rect 25228 37874 25284 37884
rect 23884 37380 23940 37390
rect 23884 36708 23940 37324
rect 24444 37266 24500 37436
rect 24444 37214 24446 37266
rect 24498 37214 24500 37266
rect 24444 37202 24500 37214
rect 24556 37604 24612 37614
rect 23884 36642 23940 36652
rect 23996 36596 24052 36606
rect 23996 36370 24052 36540
rect 24220 36596 24276 36606
rect 23996 36318 23998 36370
rect 24050 36318 24052 36370
rect 23996 36306 24052 36318
rect 24108 36484 24164 36494
rect 23884 36258 23940 36270
rect 23884 36206 23886 36258
rect 23938 36206 23940 36258
rect 23884 35810 23940 36206
rect 23884 35758 23886 35810
rect 23938 35758 23940 35810
rect 23884 35746 23940 35758
rect 23772 35074 23828 35084
rect 23548 34962 23604 34972
rect 23772 34914 23828 34926
rect 23772 34862 23774 34914
rect 23826 34862 23828 34914
rect 22652 34078 22654 34130
rect 22706 34078 22708 34130
rect 22652 34066 22708 34078
rect 22988 34524 23380 34580
rect 23548 34802 23604 34814
rect 23548 34750 23550 34802
rect 23602 34750 23604 34802
rect 23548 34580 23604 34750
rect 23772 34804 23828 34862
rect 23772 34738 23828 34748
rect 24108 34580 24164 36428
rect 23604 34524 24164 34580
rect 22316 33404 22484 33460
rect 22540 33404 22820 33460
rect 22428 33348 22484 33404
rect 22428 33292 22596 33348
rect 22204 31668 22260 33068
rect 22316 33236 22372 33246
rect 22316 32674 22372 33180
rect 22428 33122 22484 33134
rect 22428 33070 22430 33122
rect 22482 33070 22484 33122
rect 22428 32788 22484 33070
rect 22428 32722 22484 32732
rect 22316 32622 22318 32674
rect 22370 32622 22372 32674
rect 22316 32610 22372 32622
rect 22428 31780 22484 31790
rect 22428 31686 22484 31724
rect 22204 31602 22260 31612
rect 22540 31332 22596 33292
rect 22428 31276 22596 31332
rect 22428 30548 22484 31276
rect 22652 31220 22708 31230
rect 22428 30482 22484 30492
rect 22540 31108 22596 31118
rect 22092 30156 22260 30212
rect 21308 30098 21364 30110
rect 21308 30046 21310 30098
rect 21362 30046 21364 30098
rect 21308 29652 21364 30046
rect 21308 29586 21364 29596
rect 21196 29374 21198 29426
rect 21250 29374 21252 29426
rect 21196 29362 21252 29374
rect 21532 28868 21588 28878
rect 21644 28868 21700 30156
rect 21756 30146 21812 30156
rect 21980 30100 22036 30110
rect 21980 30006 22036 30044
rect 22204 29764 22260 30156
rect 22428 30210 22484 30222
rect 22428 30158 22430 30210
rect 22482 30158 22484 30210
rect 22428 29988 22484 30158
rect 22428 29922 22484 29932
rect 22092 29708 22260 29764
rect 21756 29428 21812 29438
rect 21756 29334 21812 29372
rect 21532 28866 21700 28868
rect 21532 28814 21534 28866
rect 21586 28814 21700 28866
rect 21532 28812 21700 28814
rect 21532 28802 21588 28812
rect 21980 28642 22036 28654
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21644 28532 21700 28542
rect 21980 28532 22036 28590
rect 21644 28530 22036 28532
rect 21644 28478 21646 28530
rect 21698 28478 22036 28530
rect 21644 28476 22036 28478
rect 21644 28466 21700 28476
rect 21532 28420 21588 28430
rect 21420 28418 21588 28420
rect 21420 28366 21534 28418
rect 21586 28366 21588 28418
rect 21420 28364 21588 28366
rect 21420 26964 21476 28364
rect 21532 28354 21588 28364
rect 21644 28308 21700 28318
rect 21532 28196 21588 28206
rect 21532 27858 21588 28140
rect 21644 27970 21700 28252
rect 21644 27918 21646 27970
rect 21698 27918 21700 27970
rect 21644 27906 21700 27918
rect 21532 27806 21534 27858
rect 21586 27806 21588 27858
rect 21532 27794 21588 27806
rect 21644 27188 21700 27198
rect 21756 27188 21812 28476
rect 21700 27132 21812 27188
rect 21644 27122 21700 27132
rect 21084 26852 21252 26908
rect 19964 25620 20020 25630
rect 19852 25618 20020 25620
rect 19852 25566 19966 25618
rect 20018 25566 20020 25618
rect 19852 25564 20020 25566
rect 19964 25554 20020 25564
rect 19292 25454 19294 25506
rect 19346 25454 19348 25506
rect 19292 25442 19348 25454
rect 20076 25506 20132 25518
rect 20076 25454 20078 25506
rect 20130 25454 20132 25506
rect 20076 25284 20132 25454
rect 20076 25218 20132 25228
rect 20412 25394 20468 25406
rect 20412 25342 20414 25394
rect 20466 25342 20468 25394
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19180 24558 19182 24610
rect 19234 24558 19236 24610
rect 19180 24546 19236 24558
rect 19292 24834 19348 24846
rect 20412 24836 20468 25342
rect 19292 24782 19294 24834
rect 19346 24782 19348 24834
rect 18620 24220 19236 24276
rect 18228 23772 18564 23828
rect 19068 23828 19124 23838
rect 18172 23734 18228 23772
rect 16604 23380 16660 23390
rect 16492 23378 16660 23380
rect 16492 23326 16606 23378
rect 16658 23326 16660 23378
rect 16492 23324 16660 23326
rect 16604 23314 16660 23324
rect 19068 23378 19124 23772
rect 19068 23326 19070 23378
rect 19122 23326 19124 23378
rect 19068 23314 19124 23326
rect 19180 23266 19236 24220
rect 19180 23214 19182 23266
rect 19234 23214 19236 23266
rect 19180 23202 19236 23214
rect 17612 23042 17668 23054
rect 17612 22990 17614 23042
rect 17666 22990 17668 23042
rect 16156 22932 16212 22942
rect 16044 22876 16156 22932
rect 16156 22866 16212 22876
rect 17612 22932 17668 22990
rect 17612 22866 17668 22876
rect 19068 22932 19124 22942
rect 19292 22932 19348 24782
rect 20300 24834 20468 24836
rect 20300 24782 20414 24834
rect 20466 24782 20468 24834
rect 20300 24780 20468 24782
rect 19964 24724 20020 24734
rect 19740 24052 19796 24062
rect 19740 23958 19796 23996
rect 19964 23938 20020 24668
rect 19964 23886 19966 23938
rect 20018 23886 20020 23938
rect 19964 23874 20020 23886
rect 20188 23940 20244 23950
rect 20188 23846 20244 23884
rect 20300 23938 20356 24780
rect 20412 24770 20468 24780
rect 20636 24164 20692 26852
rect 21196 26516 21252 26852
rect 20860 26404 20916 26414
rect 20860 26310 20916 26348
rect 21196 26290 21252 26460
rect 21196 26238 21198 26290
rect 21250 26238 21252 26290
rect 21196 26226 21252 26238
rect 20972 24836 21028 24846
rect 20748 24164 20804 24174
rect 20636 24162 20804 24164
rect 20636 24110 20750 24162
rect 20802 24110 20804 24162
rect 20636 24108 20804 24110
rect 20748 24098 20804 24108
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 20300 23874 20356 23886
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20972 23548 21028 24780
rect 21084 24722 21140 24734
rect 21084 24670 21086 24722
rect 21138 24670 21140 24722
rect 21084 23940 21140 24670
rect 21084 23828 21140 23884
rect 21308 23828 21364 23838
rect 21084 23826 21364 23828
rect 21084 23774 21310 23826
rect 21362 23774 21364 23826
rect 21084 23772 21364 23774
rect 21308 23762 21364 23772
rect 20972 23492 21140 23548
rect 19836 23482 20100 23492
rect 21084 23378 21140 23492
rect 21084 23326 21086 23378
rect 21138 23326 21140 23378
rect 21084 23314 21140 23326
rect 21308 23268 21364 23278
rect 21420 23268 21476 26908
rect 21980 26852 22036 26862
rect 21756 26796 21980 26852
rect 21756 26514 21812 26796
rect 21980 26758 22036 26796
rect 21756 26462 21758 26514
rect 21810 26462 21812 26514
rect 21756 26450 21812 26462
rect 21756 25506 21812 25518
rect 21756 25454 21758 25506
rect 21810 25454 21812 25506
rect 21532 25284 21588 25294
rect 21756 25284 21812 25454
rect 21588 25228 21812 25284
rect 21868 25284 21924 25294
rect 22092 25284 22148 29708
rect 22204 29428 22260 29438
rect 22204 26852 22260 29372
rect 22540 28642 22596 31052
rect 22652 30098 22708 31164
rect 22652 30046 22654 30098
rect 22706 30046 22708 30098
rect 22652 29652 22708 30046
rect 22652 29586 22708 29596
rect 22540 28590 22542 28642
rect 22594 28590 22596 28642
rect 22540 28578 22596 28590
rect 22652 29314 22708 29326
rect 22652 29262 22654 29314
rect 22706 29262 22708 29314
rect 22652 28644 22708 29262
rect 22204 26290 22260 26796
rect 22204 26238 22206 26290
rect 22258 26238 22260 26290
rect 22204 26180 22260 26238
rect 22204 26114 22260 26124
rect 21868 25282 22148 25284
rect 21868 25230 21870 25282
rect 21922 25230 22148 25282
rect 21868 25228 22148 25230
rect 22540 25394 22596 25406
rect 22540 25342 22542 25394
rect 22594 25342 22596 25394
rect 21532 25190 21588 25228
rect 21868 25218 21924 25228
rect 21532 24836 21588 24846
rect 21532 24050 21588 24780
rect 22428 24834 22484 24846
rect 22428 24782 22430 24834
rect 22482 24782 22484 24834
rect 21980 24722 22036 24734
rect 21980 24670 21982 24722
rect 22034 24670 22036 24722
rect 21980 24164 22036 24670
rect 21980 24098 22036 24108
rect 22316 24164 22372 24174
rect 21532 23998 21534 24050
rect 21586 23998 21588 24050
rect 21532 23986 21588 23998
rect 21980 23938 22036 23950
rect 21980 23886 21982 23938
rect 22034 23886 22036 23938
rect 21644 23380 21700 23390
rect 21980 23380 22036 23886
rect 22316 23938 22372 24108
rect 22316 23886 22318 23938
rect 22370 23886 22372 23938
rect 22316 23874 22372 23886
rect 22428 23492 22484 24782
rect 22540 24164 22596 25342
rect 22652 25284 22708 28588
rect 22764 26178 22820 33404
rect 22876 33124 22932 33134
rect 22876 32564 22932 33068
rect 22876 32498 22932 32508
rect 22876 31780 22932 31790
rect 22876 31108 22932 31724
rect 22876 31042 22932 31052
rect 22876 30548 22932 30558
rect 22876 27188 22932 30492
rect 22988 29876 23044 34524
rect 23548 34514 23604 34524
rect 23548 34130 23604 34142
rect 23548 34078 23550 34130
rect 23602 34078 23604 34130
rect 23212 33460 23268 33470
rect 23212 33366 23268 33404
rect 23324 33348 23380 33358
rect 23324 33254 23380 33292
rect 23548 33236 23604 34078
rect 23548 33170 23604 33180
rect 23100 33122 23156 33134
rect 23100 33070 23102 33122
rect 23154 33070 23156 33122
rect 23100 33012 23156 33070
rect 23100 32946 23156 32956
rect 23212 33124 23268 33134
rect 23212 32450 23268 33068
rect 23660 33124 23716 34524
rect 23884 34244 23940 34254
rect 23660 33058 23716 33068
rect 23772 34242 23940 34244
rect 23772 34190 23886 34242
rect 23938 34190 23940 34242
rect 23772 34188 23940 34190
rect 23772 33346 23828 34188
rect 23884 34178 23940 34188
rect 24220 34242 24276 36540
rect 24444 36596 24500 36606
rect 24332 35364 24388 35374
rect 24332 34804 24388 35308
rect 24332 34738 24388 34748
rect 24220 34190 24222 34242
rect 24274 34190 24276 34242
rect 24220 34178 24276 34190
rect 23996 34132 24052 34142
rect 23996 34038 24052 34076
rect 23772 33294 23774 33346
rect 23826 33294 23828 33346
rect 23212 32398 23214 32450
rect 23266 32398 23268 32450
rect 23212 32386 23268 32398
rect 23660 32562 23716 32574
rect 23660 32510 23662 32562
rect 23714 32510 23716 32562
rect 23212 32004 23268 32014
rect 23212 30324 23268 31948
rect 23660 31780 23716 32510
rect 23660 31714 23716 31724
rect 23772 31668 23828 33294
rect 24220 31668 24276 31678
rect 23772 31666 24276 31668
rect 23772 31614 24222 31666
rect 24274 31614 24276 31666
rect 23772 31612 24276 31614
rect 23212 30258 23268 30268
rect 23772 30996 23828 31006
rect 23100 30212 23156 30222
rect 23100 30098 23156 30156
rect 23548 30210 23604 30222
rect 23548 30158 23550 30210
rect 23602 30158 23604 30210
rect 23324 30100 23380 30110
rect 23100 30046 23102 30098
rect 23154 30046 23156 30098
rect 23100 30034 23156 30046
rect 23212 30098 23380 30100
rect 23212 30046 23326 30098
rect 23378 30046 23380 30098
rect 23212 30044 23380 30046
rect 22988 29820 23156 29876
rect 22988 28084 23044 28094
rect 22988 27990 23044 28028
rect 22876 27122 22932 27132
rect 23100 26908 23156 29820
rect 23212 28756 23268 30044
rect 23324 30034 23380 30044
rect 23548 29988 23604 30158
rect 23436 29652 23492 29662
rect 23436 29558 23492 29596
rect 23548 29316 23604 29932
rect 23772 29764 23828 30940
rect 23996 30212 24052 30222
rect 23772 29650 23828 29708
rect 23772 29598 23774 29650
rect 23826 29598 23828 29650
rect 23772 29540 23828 29598
rect 23884 30100 23940 30110
rect 23884 29652 23940 30044
rect 23996 30098 24052 30156
rect 23996 30046 23998 30098
rect 24050 30046 24052 30098
rect 23996 30034 24052 30046
rect 23996 29652 24052 29662
rect 23884 29650 24052 29652
rect 23884 29598 23998 29650
rect 24050 29598 24052 29650
rect 23884 29596 24052 29598
rect 23996 29586 24052 29596
rect 23772 29474 23828 29484
rect 24108 29428 24164 31612
rect 24220 31602 24276 31612
rect 24220 31444 24276 31454
rect 24220 31218 24276 31388
rect 24220 31166 24222 31218
rect 24274 31166 24276 31218
rect 24220 31154 24276 31166
rect 24444 30996 24500 36540
rect 24556 31890 24612 37548
rect 24668 37490 24724 37502
rect 24668 37438 24670 37490
rect 24722 37438 24724 37490
rect 24668 35700 24724 37438
rect 25340 35812 25396 37884
rect 25452 37154 25508 37166
rect 25452 37102 25454 37154
rect 25506 37102 25508 37154
rect 25452 36484 25508 37102
rect 25452 36418 25508 36428
rect 25228 35700 25284 35710
rect 24668 35698 25284 35700
rect 24668 35646 25230 35698
rect 25282 35646 25284 35698
rect 24668 35644 25284 35646
rect 25228 35634 25284 35644
rect 25340 35586 25396 35756
rect 25340 35534 25342 35586
rect 25394 35534 25396 35586
rect 25340 35522 25396 35534
rect 25452 35810 25508 35822
rect 25452 35758 25454 35810
rect 25506 35758 25508 35810
rect 25340 35140 25396 35150
rect 25228 34914 25284 34926
rect 25228 34862 25230 34914
rect 25282 34862 25284 34914
rect 24668 34018 24724 34030
rect 24668 33966 24670 34018
rect 24722 33966 24724 34018
rect 24668 33796 24724 33966
rect 24668 33730 24724 33740
rect 24780 33572 24836 33582
rect 24668 32788 24724 32798
rect 24668 32694 24724 32732
rect 24556 31838 24558 31890
rect 24610 31838 24612 31890
rect 24556 31826 24612 31838
rect 24780 31218 24836 33516
rect 25228 33460 25284 34862
rect 25340 34802 25396 35084
rect 25340 34750 25342 34802
rect 25394 34750 25396 34802
rect 25340 34738 25396 34750
rect 25452 34356 25508 35758
rect 25452 34290 25508 34300
rect 25340 34130 25396 34142
rect 25564 34132 25620 34142
rect 25340 34078 25342 34130
rect 25394 34078 25396 34130
rect 25340 33684 25396 34078
rect 25340 33618 25396 33628
rect 25452 34130 25620 34132
rect 25452 34078 25566 34130
rect 25618 34078 25620 34130
rect 25452 34076 25620 34078
rect 25228 33394 25284 33404
rect 25116 33236 25172 33246
rect 24892 31780 24948 31790
rect 25116 31780 25172 33180
rect 25452 32788 25508 34076
rect 25564 34066 25620 34076
rect 24892 31778 25172 31780
rect 24892 31726 24894 31778
rect 24946 31726 25172 31778
rect 24892 31724 25172 31726
rect 25340 32564 25396 32574
rect 24892 31714 24948 31724
rect 25228 31668 25284 31678
rect 24780 31166 24782 31218
rect 24834 31166 24836 31218
rect 24780 31154 24836 31166
rect 25004 31666 25284 31668
rect 25004 31614 25230 31666
rect 25282 31614 25284 31666
rect 25004 31612 25284 31614
rect 24444 30940 24836 30996
rect 24668 30436 24724 30446
rect 24332 30324 24388 30334
rect 24332 30098 24388 30268
rect 24332 30046 24334 30098
rect 24386 30046 24388 30098
rect 24332 30034 24388 30046
rect 24220 29764 24276 29774
rect 24220 29650 24276 29708
rect 24220 29598 24222 29650
rect 24274 29598 24276 29650
rect 24220 29586 24276 29598
rect 23548 29250 23604 29260
rect 23996 29372 24164 29428
rect 24332 29426 24388 29438
rect 24332 29374 24334 29426
rect 24386 29374 24388 29426
rect 23212 28690 23268 28700
rect 23324 28644 23380 28654
rect 23324 28550 23380 28588
rect 23436 28532 23492 28542
rect 23436 28438 23492 28476
rect 23772 27188 23828 27198
rect 23772 27094 23828 27132
rect 23996 26908 24052 29372
rect 24332 29204 24388 29374
rect 24220 28530 24276 28542
rect 24220 28478 24222 28530
rect 24274 28478 24276 28530
rect 24220 28084 24276 28478
rect 24332 28420 24388 29148
rect 24556 28756 24612 28766
rect 24556 28662 24612 28700
rect 24668 28642 24724 30380
rect 24668 28590 24670 28642
rect 24722 28590 24724 28642
rect 24668 28532 24724 28590
rect 24332 28354 24388 28364
rect 24556 28476 24724 28532
rect 24220 28018 24276 28028
rect 24220 27188 24276 27198
rect 24220 27074 24276 27132
rect 24220 27022 24222 27074
rect 24274 27022 24276 27074
rect 24220 27010 24276 27022
rect 24444 27074 24500 27086
rect 24444 27022 24446 27074
rect 24498 27022 24500 27074
rect 23100 26852 23380 26908
rect 23996 26852 24276 26908
rect 22764 26126 22766 26178
rect 22818 26126 22820 26178
rect 22764 25396 22820 26126
rect 23212 26180 23268 26190
rect 23100 25844 23156 25854
rect 22764 25330 22820 25340
rect 22988 25788 23100 25844
rect 22652 25218 22708 25228
rect 22988 24946 23044 25788
rect 23100 25778 23156 25788
rect 23212 25172 23268 26124
rect 23212 25106 23268 25116
rect 22988 24894 22990 24946
rect 23042 24894 23044 24946
rect 22988 24882 23044 24894
rect 23324 24836 23380 26852
rect 23660 26068 23716 26078
rect 22540 24098 22596 24108
rect 23100 24780 23324 24836
rect 22428 23426 22484 23436
rect 21644 23378 22036 23380
rect 21644 23326 21646 23378
rect 21698 23326 22036 23378
rect 21644 23324 22036 23326
rect 21644 23314 21700 23324
rect 21364 23212 21476 23268
rect 21980 23268 22036 23324
rect 22988 23380 23044 23390
rect 23100 23380 23156 24780
rect 23324 24770 23380 24780
rect 23436 25732 23492 25742
rect 23436 24050 23492 25676
rect 23660 25506 23716 26012
rect 24220 25844 24276 26852
rect 24220 25778 24276 25788
rect 24444 25732 24500 27022
rect 24444 25666 24500 25676
rect 23660 25454 23662 25506
rect 23714 25454 23716 25506
rect 23660 25442 23716 25454
rect 23548 25396 23604 25406
rect 23548 25302 23604 25340
rect 24444 25172 24500 25182
rect 23436 23998 23438 24050
rect 23490 23998 23492 24050
rect 23436 23986 23492 23998
rect 23772 24948 23828 24958
rect 23772 24052 23828 24892
rect 24220 24836 24276 24846
rect 24220 24742 24276 24780
rect 24444 24722 24500 25116
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 24220 24052 24276 24062
rect 23772 24050 24276 24052
rect 23772 23998 24222 24050
rect 24274 23998 24276 24050
rect 23772 23996 24276 23998
rect 23772 23938 23828 23996
rect 24220 23986 24276 23996
rect 24444 24052 24500 24670
rect 24444 23986 24500 23996
rect 23772 23886 23774 23938
rect 23826 23886 23828 23938
rect 23772 23874 23828 23886
rect 24556 23828 24612 28476
rect 24668 27748 24724 27758
rect 24668 27654 24724 27692
rect 24668 27300 24724 27310
rect 24780 27300 24836 30940
rect 25004 30212 25060 31612
rect 25228 31602 25284 31612
rect 25004 30118 25060 30156
rect 25116 30996 25172 31006
rect 25116 30324 25172 30940
rect 25340 30882 25396 32508
rect 25340 30830 25342 30882
rect 25394 30830 25396 30882
rect 25340 30818 25396 30830
rect 25452 30660 25508 32732
rect 25564 33346 25620 33358
rect 25564 33294 25566 33346
rect 25618 33294 25620 33346
rect 25564 32004 25620 33294
rect 25564 31938 25620 31948
rect 25116 30210 25172 30268
rect 25116 30158 25118 30210
rect 25170 30158 25172 30210
rect 25116 30146 25172 30158
rect 25340 30604 25508 30660
rect 25228 30098 25284 30110
rect 25228 30046 25230 30098
rect 25282 30046 25284 30098
rect 25228 29988 25284 30046
rect 25228 29922 25284 29932
rect 25116 28644 25172 28654
rect 25116 28550 25172 28588
rect 24668 27298 24836 27300
rect 24668 27246 24670 27298
rect 24722 27246 24836 27298
rect 24668 27244 24836 27246
rect 24668 27234 24724 27244
rect 25228 27076 25284 27086
rect 25228 26982 25284 27020
rect 25228 26628 25284 26638
rect 25228 26292 25284 26572
rect 25340 26404 25396 30604
rect 25676 30436 25732 40124
rect 26348 40114 26404 40124
rect 25788 39844 25844 39854
rect 26124 39844 26180 39854
rect 25844 39788 26068 39844
rect 25788 39778 25844 39788
rect 25900 39508 25956 39518
rect 25788 39506 25956 39508
rect 25788 39454 25902 39506
rect 25954 39454 25956 39506
rect 25788 39452 25956 39454
rect 25788 38610 25844 39452
rect 25900 39442 25956 39452
rect 26012 38834 26068 39788
rect 26012 38782 26014 38834
rect 26066 38782 26068 38834
rect 26012 38770 26068 38782
rect 26124 38668 26180 39788
rect 26348 39508 26404 39518
rect 26236 38948 26292 38958
rect 26236 38854 26292 38892
rect 26348 38668 26404 39452
rect 25788 38558 25790 38610
rect 25842 38558 25844 38610
rect 25788 37604 25844 38558
rect 25788 37538 25844 37548
rect 25900 38612 26180 38668
rect 26236 38612 26404 38668
rect 25788 37380 25844 37390
rect 25788 37286 25844 37324
rect 25788 37044 25844 37054
rect 25788 36482 25844 36988
rect 25788 36430 25790 36482
rect 25842 36430 25844 36482
rect 25788 36418 25844 36430
rect 25900 36596 25956 38612
rect 26124 38052 26180 38062
rect 26124 37958 26180 37996
rect 26124 37492 26180 37502
rect 26124 37378 26180 37436
rect 26124 37326 26126 37378
rect 26178 37326 26180 37378
rect 26124 37314 26180 37326
rect 25788 35476 25844 35486
rect 25788 31220 25844 35420
rect 25900 34802 25956 36540
rect 25900 34750 25902 34802
rect 25954 34750 25956 34802
rect 25900 34242 25956 34750
rect 26012 36482 26068 36494
rect 26012 36430 26014 36482
rect 26066 36430 26068 36482
rect 26012 34804 26068 36430
rect 26012 34738 26068 34748
rect 26236 35028 26292 38612
rect 26460 37492 26516 44380
rect 26908 44324 26964 44334
rect 27132 44324 27188 48190
rect 27356 46676 27412 48302
rect 27468 47458 27524 48524
rect 27468 47406 27470 47458
rect 27522 47406 27524 47458
rect 27468 47394 27524 47406
rect 27580 47012 27636 49420
rect 27692 47460 27748 49534
rect 27916 49028 27972 49038
rect 27916 48934 27972 48972
rect 27692 47394 27748 47404
rect 27804 48692 27860 48702
rect 27580 46946 27636 46956
rect 27804 47346 27860 48636
rect 28028 48580 28084 51884
rect 28252 51268 28308 51278
rect 28252 51174 28308 51212
rect 28364 51044 28420 55804
rect 30044 55468 30100 56142
rect 30268 56082 30324 56364
rect 31724 56308 31780 56318
rect 32060 56308 32116 59200
rect 34300 56308 34356 59200
rect 36540 56308 36596 59200
rect 38780 56642 38836 59200
rect 38780 56590 38782 56642
rect 38834 56590 38836 56642
rect 38780 56578 38836 56590
rect 39340 56642 39396 56654
rect 39340 56590 39342 56642
rect 39394 56590 39396 56642
rect 31724 56306 32340 56308
rect 31724 56254 31726 56306
rect 31778 56254 32340 56306
rect 31724 56252 32340 56254
rect 31724 56242 31780 56252
rect 32284 56194 32340 56252
rect 34300 56306 34580 56308
rect 34300 56254 34302 56306
rect 34354 56254 34580 56306
rect 34300 56252 34580 56254
rect 34300 56242 34356 56252
rect 32284 56142 32286 56194
rect 32338 56142 32340 56194
rect 32284 56130 32340 56142
rect 32620 56194 32676 56206
rect 32620 56142 32622 56194
rect 32674 56142 32676 56194
rect 30268 56030 30270 56082
rect 30322 56030 30324 56082
rect 30268 56018 30324 56030
rect 29372 55412 30100 55468
rect 29260 55300 29316 55310
rect 29260 55206 29316 55244
rect 29148 54628 29204 54638
rect 29204 54572 29316 54628
rect 29148 54534 29204 54572
rect 28812 54516 28868 54526
rect 28812 54422 28868 54460
rect 29260 53956 29316 54572
rect 29372 54180 29428 55412
rect 32060 55410 32116 55422
rect 32060 55358 32062 55410
rect 32114 55358 32116 55410
rect 29932 55186 29988 55198
rect 29932 55134 29934 55186
rect 29986 55134 29988 55186
rect 29484 54740 29540 54750
rect 29484 54738 29876 54740
rect 29484 54686 29486 54738
rect 29538 54686 29876 54738
rect 29484 54684 29876 54686
rect 29484 54674 29540 54684
rect 29820 54514 29876 54684
rect 29932 54738 29988 55134
rect 29932 54686 29934 54738
rect 29986 54686 29988 54738
rect 29932 54674 29988 54686
rect 31836 54628 31892 54638
rect 29820 54462 29822 54514
rect 29874 54462 29876 54514
rect 29372 54124 29652 54180
rect 29260 53842 29316 53900
rect 29260 53790 29262 53842
rect 29314 53790 29316 53842
rect 29260 53778 29316 53790
rect 29148 53508 29204 53518
rect 29148 53170 29204 53452
rect 29148 53118 29150 53170
rect 29202 53118 29204 53170
rect 29148 53106 29204 53118
rect 29596 53058 29652 54124
rect 29596 53006 29598 53058
rect 29650 53006 29652 53058
rect 29596 52994 29652 53006
rect 29820 53060 29876 54462
rect 30044 54516 30100 54526
rect 30044 54422 30100 54460
rect 30604 54516 30660 54526
rect 30604 54514 31780 54516
rect 30604 54462 30606 54514
rect 30658 54462 31780 54514
rect 30604 54460 31780 54462
rect 30604 54450 30660 54460
rect 31724 54402 31780 54460
rect 31724 54350 31726 54402
rect 31778 54350 31780 54402
rect 31724 54338 31780 54350
rect 30380 54290 30436 54302
rect 30380 54238 30382 54290
rect 30434 54238 30436 54290
rect 30380 53844 30436 54238
rect 30156 53508 30212 53518
rect 29932 53060 29988 53070
rect 29820 53004 29932 53060
rect 29932 52966 29988 53004
rect 30156 53058 30212 53452
rect 30156 53006 30158 53058
rect 30210 53006 30212 53058
rect 30156 52994 30212 53006
rect 30380 52946 30436 53788
rect 31836 53172 31892 54572
rect 32060 54290 32116 55358
rect 32620 55298 32676 56142
rect 34524 56194 34580 56252
rect 36540 56306 36820 56308
rect 36540 56254 36542 56306
rect 36594 56254 36820 56306
rect 36540 56252 36820 56254
rect 36540 56242 36596 56252
rect 34524 56142 34526 56194
rect 34578 56142 34580 56194
rect 34524 56130 34580 56142
rect 34860 56194 34916 56206
rect 34860 56142 34862 56194
rect 34914 56142 34916 56194
rect 32620 55246 32622 55298
rect 32674 55246 32676 55298
rect 32620 55234 32676 55246
rect 33180 55300 33236 55310
rect 32508 55076 32564 55086
rect 32508 54738 32564 55020
rect 32620 55076 32676 55086
rect 33180 55076 33236 55244
rect 33628 55298 33684 55310
rect 33628 55246 33630 55298
rect 33682 55246 33684 55298
rect 33628 55076 33684 55246
rect 32620 55074 32788 55076
rect 32620 55022 32622 55074
rect 32674 55022 32788 55074
rect 32620 55020 32788 55022
rect 32620 55010 32676 55020
rect 32508 54686 32510 54738
rect 32562 54686 32564 54738
rect 32508 54628 32564 54686
rect 32508 54562 32564 54572
rect 32060 54238 32062 54290
rect 32114 54238 32116 54290
rect 32060 53732 32116 54238
rect 32060 53666 32116 53676
rect 32620 53620 32676 53630
rect 32620 53526 32676 53564
rect 31948 53172 32004 53182
rect 31836 53170 32004 53172
rect 31836 53118 31950 53170
rect 32002 53118 32004 53170
rect 31836 53116 32004 53118
rect 31948 53106 32004 53116
rect 32172 53060 32228 53070
rect 32228 53004 32340 53060
rect 32172 52966 32228 53004
rect 30380 52894 30382 52946
rect 30434 52894 30436 52946
rect 30380 52882 30436 52894
rect 30716 52948 30772 52958
rect 30716 52854 30772 52892
rect 31836 52948 31892 52958
rect 30044 52834 30100 52846
rect 30044 52782 30046 52834
rect 30098 52782 30100 52834
rect 29484 52722 29540 52734
rect 29484 52670 29486 52722
rect 29538 52670 29540 52722
rect 29372 52164 29428 52174
rect 29372 52070 29428 52108
rect 29484 52052 29540 52670
rect 30044 52276 30100 52782
rect 31836 52834 31892 52892
rect 31836 52782 31838 52834
rect 31890 52782 31892 52834
rect 31836 52770 31892 52782
rect 30156 52276 30212 52286
rect 30044 52274 30212 52276
rect 30044 52222 30158 52274
rect 30210 52222 30212 52274
rect 30044 52220 30212 52222
rect 30156 52210 30212 52220
rect 32284 52274 32340 53004
rect 32732 52500 32788 55020
rect 33180 55074 33684 55076
rect 33180 55022 33182 55074
rect 33234 55022 33684 55074
rect 33180 55020 33684 55022
rect 33180 55010 33236 55020
rect 33404 54628 33460 54638
rect 33628 54628 33684 55020
rect 34300 55186 34356 55198
rect 34300 55134 34302 55186
rect 34354 55134 34356 55186
rect 33964 54740 34020 54750
rect 34300 54740 34356 55134
rect 33964 54738 34356 54740
rect 33964 54686 33966 54738
rect 34018 54686 34356 54738
rect 33964 54684 34356 54686
rect 33964 54674 34020 54684
rect 33404 54534 33460 54572
rect 33516 54572 33628 54628
rect 33180 54514 33236 54526
rect 33180 54462 33182 54514
rect 33234 54462 33236 54514
rect 33068 53730 33124 53742
rect 33068 53678 33070 53730
rect 33122 53678 33124 53730
rect 33068 53620 33124 53678
rect 33068 53554 33124 53564
rect 33180 53172 33236 54462
rect 33292 53844 33348 53854
rect 33292 53618 33348 53788
rect 33292 53566 33294 53618
rect 33346 53566 33348 53618
rect 33292 53554 33348 53566
rect 33068 53060 33124 53070
rect 33180 53060 33236 53116
rect 33068 53058 33236 53060
rect 33068 53006 33070 53058
rect 33122 53006 33236 53058
rect 33068 53004 33236 53006
rect 33068 52994 33124 53004
rect 32284 52222 32286 52274
rect 32338 52222 32340 52274
rect 32284 52210 32340 52222
rect 32620 52444 32788 52500
rect 33292 52946 33348 52958
rect 33292 52894 33294 52946
rect 33346 52894 33348 52946
rect 29484 51986 29540 51996
rect 28252 50988 28420 51044
rect 32620 51268 32676 52444
rect 32732 52276 32788 52286
rect 33292 52276 33348 52894
rect 32788 52220 33348 52276
rect 32732 52182 32788 52220
rect 33404 52164 33460 52174
rect 33516 52164 33572 54572
rect 33628 54562 33684 54572
rect 33852 54516 33908 54526
rect 33628 54290 33684 54302
rect 33628 54238 33630 54290
rect 33682 54238 33684 54290
rect 33628 53844 33684 54238
rect 33628 52722 33684 53788
rect 33852 53620 33908 54460
rect 33964 54514 34020 54526
rect 33964 54462 33966 54514
rect 34018 54462 34020 54514
rect 33964 54404 34020 54462
rect 34860 54514 34916 56142
rect 36764 56194 36820 56252
rect 39340 56306 39396 56590
rect 39340 56254 39342 56306
rect 39394 56254 39396 56306
rect 39340 56242 39396 56254
rect 40124 56642 40180 56654
rect 40124 56590 40126 56642
rect 40178 56590 40180 56642
rect 36764 56142 36766 56194
rect 36818 56142 36820 56194
rect 36764 56130 36820 56142
rect 37100 56194 37156 56206
rect 37100 56142 37102 56194
rect 37154 56142 37156 56194
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 36428 55410 36484 55422
rect 36428 55358 36430 55410
rect 36482 55358 36484 55410
rect 36092 54740 36148 54750
rect 36092 54628 36148 54684
rect 36204 54628 36260 54638
rect 36092 54626 36260 54628
rect 36092 54574 36206 54626
rect 36258 54574 36260 54626
rect 36092 54572 36260 54574
rect 36204 54562 36260 54572
rect 34860 54462 34862 54514
rect 34914 54462 34916 54514
rect 34860 54450 34916 54462
rect 33964 54338 34020 54348
rect 34748 54402 34804 54414
rect 34748 54350 34750 54402
rect 34802 54350 34804 54402
rect 33852 53554 33908 53564
rect 34636 53620 34692 53630
rect 33852 53172 33908 53182
rect 33852 53170 34132 53172
rect 33852 53118 33854 53170
rect 33906 53118 34132 53170
rect 33852 53116 34132 53118
rect 33852 53106 33908 53116
rect 33852 52948 33908 52958
rect 33852 52854 33908 52892
rect 33628 52670 33630 52722
rect 33682 52670 33684 52722
rect 33628 52658 33684 52670
rect 34076 52274 34132 53116
rect 34076 52222 34078 52274
rect 34130 52222 34132 52274
rect 34076 52210 34132 52222
rect 28028 48514 28084 48524
rect 28140 49140 28196 49150
rect 28140 48356 28196 49084
rect 27804 47294 27806 47346
rect 27858 47294 27860 47346
rect 27356 46620 27524 46676
rect 27356 45780 27412 45790
rect 27356 45686 27412 45724
rect 27468 45332 27524 46620
rect 27580 45332 27636 45342
rect 27468 45330 27636 45332
rect 27468 45278 27582 45330
rect 27634 45278 27636 45330
rect 27468 45276 27636 45278
rect 27580 45266 27636 45276
rect 27804 44434 27860 47294
rect 27804 44382 27806 44434
rect 27858 44382 27860 44434
rect 27804 44370 27860 44382
rect 28028 48300 28196 48356
rect 26908 44322 27188 44324
rect 26908 44270 26910 44322
rect 26962 44270 27188 44322
rect 26908 44268 27188 44270
rect 26572 44212 26628 44250
rect 26572 44146 26628 44156
rect 26796 44210 26852 44222
rect 26796 44158 26798 44210
rect 26850 44158 26852 44210
rect 26572 43988 26628 43998
rect 26796 43988 26852 44158
rect 26628 43932 26852 43988
rect 26572 43922 26628 43932
rect 26572 43540 26628 43550
rect 26684 43540 26740 43550
rect 26572 43538 26684 43540
rect 26572 43486 26574 43538
rect 26626 43486 26684 43538
rect 26572 43484 26684 43486
rect 26572 43474 26628 43484
rect 26684 43474 26740 43484
rect 26908 42084 26964 44268
rect 27132 43650 27188 43662
rect 27132 43598 27134 43650
rect 27186 43598 27188 43650
rect 27132 42980 27188 43598
rect 27244 43540 27300 43550
rect 27300 43484 27412 43540
rect 27244 43474 27300 43484
rect 27132 42914 27188 42924
rect 27020 42754 27076 42766
rect 27020 42702 27022 42754
rect 27074 42702 27076 42754
rect 27020 42308 27076 42702
rect 27020 42242 27076 42252
rect 26908 42028 27076 42084
rect 26572 41972 26628 41982
rect 26572 41878 26628 41916
rect 26908 41858 26964 41870
rect 26908 41806 26910 41858
rect 26962 41806 26964 41858
rect 26908 41412 26964 41806
rect 26908 41346 26964 41356
rect 26796 41076 26852 41086
rect 26684 40964 26740 40974
rect 26684 40626 26740 40908
rect 26684 40574 26686 40626
rect 26738 40574 26740 40626
rect 26684 40562 26740 40574
rect 26796 40404 26852 41020
rect 26684 40348 26852 40404
rect 26908 40404 26964 40414
rect 26684 39730 26740 40348
rect 26908 40292 26964 40348
rect 26684 39678 26686 39730
rect 26738 39678 26740 39730
rect 26684 39666 26740 39678
rect 26796 40236 26964 40292
rect 26796 38946 26852 40236
rect 27020 40180 27076 42028
rect 26908 40124 27076 40180
rect 27132 41410 27188 41422
rect 27132 41358 27134 41410
rect 27186 41358 27188 41410
rect 27132 40626 27188 41358
rect 27132 40574 27134 40626
rect 27186 40574 27188 40626
rect 26908 39172 26964 40124
rect 27020 39618 27076 39630
rect 27020 39566 27022 39618
rect 27074 39566 27076 39618
rect 27020 39396 27076 39566
rect 27020 39330 27076 39340
rect 26908 39116 27076 39172
rect 26796 38894 26798 38946
rect 26850 38894 26852 38946
rect 26572 38724 26628 38762
rect 26572 38658 26628 38668
rect 26796 38388 26852 38894
rect 26908 38836 26964 38846
rect 26908 38742 26964 38780
rect 26796 38332 26964 38388
rect 26684 37940 26740 37950
rect 26908 37940 26964 38332
rect 27020 38162 27076 39116
rect 27132 38834 27188 40574
rect 27244 40962 27300 40974
rect 27244 40910 27246 40962
rect 27298 40910 27300 40962
rect 27244 40404 27300 40910
rect 27244 40338 27300 40348
rect 27132 38782 27134 38834
rect 27186 38782 27188 38834
rect 27132 38770 27188 38782
rect 27356 38668 27412 43484
rect 27804 42644 27860 42654
rect 27580 41858 27636 41870
rect 27580 41806 27582 41858
rect 27634 41806 27636 41858
rect 27580 41412 27636 41806
rect 27580 41346 27636 41356
rect 27804 41300 27860 42588
rect 28028 41410 28084 48300
rect 28252 47570 28308 50988
rect 30268 50820 30324 50830
rect 30268 50596 30324 50764
rect 30268 50594 30548 50596
rect 30268 50542 30270 50594
rect 30322 50542 30548 50594
rect 30268 50540 30548 50542
rect 30268 50530 30324 50540
rect 29260 49698 29316 49710
rect 29260 49646 29262 49698
rect 29314 49646 29316 49698
rect 28588 49364 28644 49374
rect 28588 48132 28644 49308
rect 29260 48916 29316 49646
rect 29596 49140 29652 49150
rect 29260 48850 29316 48860
rect 29484 49138 29652 49140
rect 29484 49086 29598 49138
rect 29650 49086 29652 49138
rect 29484 49084 29652 49086
rect 28588 48066 28644 48076
rect 28700 48692 28756 48702
rect 28700 48242 28756 48636
rect 28700 48190 28702 48242
rect 28754 48190 28756 48242
rect 28252 47518 28254 47570
rect 28306 47518 28308 47570
rect 28252 47506 28308 47518
rect 28476 47572 28532 47582
rect 28140 44436 28196 44446
rect 28140 44322 28196 44380
rect 28140 44270 28142 44322
rect 28194 44270 28196 44322
rect 28140 44258 28196 44270
rect 28476 43708 28532 47516
rect 28700 47572 28756 48190
rect 29036 48244 29092 48254
rect 29036 48150 29092 48188
rect 28700 47506 28756 47516
rect 29148 47346 29204 47358
rect 29148 47294 29150 47346
rect 29202 47294 29204 47346
rect 28812 45668 28868 45678
rect 28140 43652 28532 43708
rect 28700 45218 28756 45230
rect 28700 45166 28702 45218
rect 28754 45166 28756 45218
rect 28140 42420 28196 43652
rect 28588 43540 28644 43550
rect 28364 43538 28644 43540
rect 28364 43486 28590 43538
rect 28642 43486 28644 43538
rect 28364 43484 28644 43486
rect 28252 43428 28308 43438
rect 28252 42866 28308 43372
rect 28364 42978 28420 43484
rect 28588 43474 28644 43484
rect 28364 42926 28366 42978
rect 28418 42926 28420 42978
rect 28364 42914 28420 42926
rect 28252 42814 28254 42866
rect 28306 42814 28308 42866
rect 28252 42802 28308 42814
rect 28476 42756 28532 42766
rect 28140 42364 28308 42420
rect 28028 41358 28030 41410
rect 28082 41358 28084 41410
rect 28028 41346 28084 41358
rect 27692 41298 27860 41300
rect 27692 41246 27806 41298
rect 27858 41246 27860 41298
rect 27692 41244 27860 41246
rect 27580 41188 27636 41198
rect 27580 39058 27636 41132
rect 27692 40068 27748 41244
rect 27804 41234 27860 41244
rect 28140 41300 28196 41310
rect 28140 41206 28196 41244
rect 28252 40404 28308 42364
rect 28476 40964 28532 42700
rect 28588 42196 28644 42206
rect 28588 42082 28644 42140
rect 28588 42030 28590 42082
rect 28642 42030 28644 42082
rect 28588 42018 28644 42030
rect 28700 41972 28756 45166
rect 28700 41906 28756 41916
rect 28588 41524 28644 41534
rect 28588 41298 28644 41468
rect 28588 41246 28590 41298
rect 28642 41246 28644 41298
rect 28588 41234 28644 41246
rect 28476 40898 28532 40908
rect 28252 40310 28308 40348
rect 28812 40402 28868 45612
rect 29148 45220 29204 47294
rect 29372 45890 29428 45902
rect 29372 45838 29374 45890
rect 29426 45838 29428 45890
rect 29148 45154 29204 45164
rect 29260 45778 29316 45790
rect 29260 45726 29262 45778
rect 29314 45726 29316 45778
rect 29148 44436 29204 44446
rect 29148 44322 29204 44380
rect 29148 44270 29150 44322
rect 29202 44270 29204 44322
rect 29148 44258 29204 44270
rect 29148 43652 29204 43662
rect 29148 43558 29204 43596
rect 29260 42194 29316 45726
rect 29372 45332 29428 45838
rect 29484 45892 29540 49084
rect 29596 49074 29652 49084
rect 30492 48466 30548 50540
rect 30604 50370 30660 50382
rect 30604 50318 30606 50370
rect 30658 50318 30660 50370
rect 30604 49140 30660 50318
rect 32396 50370 32452 50382
rect 32396 50318 32398 50370
rect 32450 50318 32452 50370
rect 32396 50036 32452 50318
rect 32508 50036 32564 50046
rect 32172 49980 32508 50036
rect 32172 49810 32228 49980
rect 32172 49758 32174 49810
rect 32226 49758 32228 49810
rect 32172 49746 32228 49758
rect 30604 49074 30660 49084
rect 31388 49698 31444 49710
rect 31388 49646 31390 49698
rect 31442 49646 31444 49698
rect 30492 48414 30494 48466
rect 30546 48414 30548 48466
rect 30492 48402 30548 48414
rect 31388 48466 31444 49646
rect 32060 49140 32116 49150
rect 31724 48916 31780 48926
rect 31388 48414 31390 48466
rect 31442 48414 31444 48466
rect 31388 48402 31444 48414
rect 31612 48914 31780 48916
rect 31612 48862 31726 48914
rect 31778 48862 31780 48914
rect 31612 48860 31780 48862
rect 29820 48356 29876 48366
rect 29820 48262 29876 48300
rect 30828 48354 30884 48366
rect 30828 48302 30830 48354
rect 30882 48302 30884 48354
rect 30828 48244 30884 48302
rect 31164 48244 31220 48254
rect 30828 48242 31220 48244
rect 30828 48190 31166 48242
rect 31218 48190 31220 48242
rect 30828 48188 31220 48190
rect 30268 47908 30324 47918
rect 29484 45826 29540 45836
rect 29596 47458 29652 47470
rect 29596 47406 29598 47458
rect 29650 47406 29652 47458
rect 29372 45266 29428 45276
rect 29596 43762 29652 47406
rect 30156 47012 30212 47022
rect 30156 46786 30212 46956
rect 30268 46900 30324 47852
rect 31164 47684 31220 48188
rect 31500 48244 31556 48254
rect 31500 48150 31556 48188
rect 31612 48020 31668 48860
rect 31724 48850 31780 48860
rect 32060 48916 32116 49084
rect 32508 49026 32564 49980
rect 32508 48974 32510 49026
rect 32562 48974 32564 49026
rect 32508 48962 32564 48974
rect 32060 48850 32116 48860
rect 31836 48804 31892 48814
rect 31724 48356 31780 48366
rect 31836 48356 31892 48748
rect 31724 48354 31892 48356
rect 31724 48302 31726 48354
rect 31778 48302 31892 48354
rect 31724 48300 31892 48302
rect 31724 48290 31780 48300
rect 32172 48244 32228 48254
rect 31612 47954 31668 47964
rect 31724 48132 31780 48142
rect 31164 47618 31220 47628
rect 30940 47572 30996 47582
rect 30940 47458 30996 47516
rect 30940 47406 30942 47458
rect 30994 47406 30996 47458
rect 30940 47394 30996 47406
rect 31276 47460 31332 47470
rect 31276 47366 31332 47404
rect 30268 46834 30324 46844
rect 31612 47124 31668 47134
rect 30156 46734 30158 46786
rect 30210 46734 30212 46786
rect 30156 46722 30212 46734
rect 30044 46228 30100 46238
rect 29596 43710 29598 43762
rect 29650 43710 29652 43762
rect 29596 43698 29652 43710
rect 29820 45106 29876 45118
rect 29820 45054 29822 45106
rect 29874 45054 29876 45106
rect 29820 44660 29876 45054
rect 29820 43708 29876 44604
rect 29932 44548 29988 44558
rect 29932 44454 29988 44492
rect 29260 42142 29262 42194
rect 29314 42142 29316 42194
rect 29260 42130 29316 42142
rect 29708 43652 29876 43708
rect 29708 41970 29764 43652
rect 29820 42756 29876 42766
rect 29820 42662 29876 42700
rect 29932 42754 29988 42766
rect 29932 42702 29934 42754
rect 29986 42702 29988 42754
rect 29932 42308 29988 42702
rect 29708 41918 29710 41970
rect 29762 41918 29764 41970
rect 29708 41906 29764 41918
rect 29820 42252 29988 42308
rect 29820 41636 29876 42252
rect 30044 42196 30100 46172
rect 30940 45890 30996 45902
rect 30940 45838 30942 45890
rect 30994 45838 30996 45890
rect 30380 44994 30436 45006
rect 30380 44942 30382 44994
rect 30434 44942 30436 44994
rect 30380 44436 30436 44942
rect 30940 44548 30996 45838
rect 30940 44482 30996 44492
rect 30380 44370 30436 44380
rect 30828 44322 30884 44334
rect 30828 44270 30830 44322
rect 30882 44270 30884 44322
rect 30604 44210 30660 44222
rect 30604 44158 30606 44210
rect 30658 44158 30660 44210
rect 30604 43988 30660 44158
rect 30604 43922 30660 43932
rect 28812 40350 28814 40402
rect 28866 40350 28868 40402
rect 28812 40338 28868 40350
rect 28924 41580 29876 41636
rect 29932 42140 30100 42196
rect 30268 43540 30324 43550
rect 27692 40002 27748 40012
rect 27804 40292 27860 40302
rect 27580 39006 27582 39058
rect 27634 39006 27636 39058
rect 27580 38994 27636 39006
rect 27804 39618 27860 40236
rect 27804 39566 27806 39618
rect 27858 39566 27860 39618
rect 27020 38110 27022 38162
rect 27074 38110 27076 38162
rect 27020 38098 27076 38110
rect 27244 38612 27412 38668
rect 27468 38948 27524 38958
rect 27468 38668 27524 38892
rect 27804 38724 27860 39566
rect 27916 40180 27972 40190
rect 28924 40180 28980 41580
rect 29372 41412 29428 41422
rect 29148 41300 29204 41310
rect 29148 41186 29204 41244
rect 29148 41134 29150 41186
rect 29202 41134 29204 41186
rect 29148 41122 29204 41134
rect 29372 41186 29428 41356
rect 29372 41134 29374 41186
rect 29426 41134 29428 41186
rect 27916 38948 27972 40124
rect 28700 40124 28980 40180
rect 29372 40852 29428 41134
rect 28588 39844 28644 39854
rect 28028 39620 28084 39630
rect 28252 39620 28308 39630
rect 28084 39564 28196 39620
rect 28028 39526 28084 39564
rect 28028 38948 28084 38958
rect 27916 38946 28084 38948
rect 27916 38894 28030 38946
rect 28082 38894 28084 38946
rect 27916 38892 28084 38894
rect 28140 38948 28196 39564
rect 28252 39618 28532 39620
rect 28252 39566 28254 39618
rect 28306 39566 28532 39618
rect 28252 39564 28532 39566
rect 28252 39554 28308 39564
rect 28140 38892 28420 38948
rect 28028 38882 28084 38892
rect 28364 38834 28420 38892
rect 28364 38782 28366 38834
rect 28418 38782 28420 38834
rect 28364 38770 28420 38782
rect 28140 38724 28196 38734
rect 27804 38722 28196 38724
rect 27804 38670 28142 38722
rect 28194 38670 28196 38722
rect 27804 38668 28196 38670
rect 27468 38612 27636 38668
rect 26684 37846 26740 37884
rect 26796 37884 26964 37940
rect 26684 37492 26740 37502
rect 26460 37490 26740 37492
rect 26460 37438 26686 37490
rect 26738 37438 26740 37490
rect 26460 37436 26740 37438
rect 26684 37426 26740 37436
rect 26460 37268 26516 37278
rect 26460 37174 26516 37212
rect 26684 35588 26740 35598
rect 26684 35364 26740 35532
rect 26684 35298 26740 35308
rect 26236 34690 26292 34972
rect 26796 35026 26852 37884
rect 26908 37604 26964 37614
rect 26908 37268 26964 37548
rect 26908 37202 26964 37212
rect 27132 37044 27188 37054
rect 27244 37044 27300 38612
rect 27132 37042 27300 37044
rect 27132 36990 27134 37042
rect 27186 36990 27300 37042
rect 27132 36988 27300 36990
rect 27132 36978 27188 36988
rect 27020 35924 27076 35934
rect 26908 35812 26964 35822
rect 26908 35364 26964 35756
rect 26908 35298 26964 35308
rect 26796 34974 26798 35026
rect 26850 34974 26852 35026
rect 26796 34962 26852 34974
rect 26236 34638 26238 34690
rect 26290 34638 26292 34690
rect 26236 34626 26292 34638
rect 26572 34914 26628 34926
rect 26572 34862 26574 34914
rect 26626 34862 26628 34914
rect 25900 34190 25902 34242
rect 25954 34190 25956 34242
rect 25900 34178 25956 34190
rect 26236 34244 26292 34254
rect 26236 34130 26292 34188
rect 26236 34078 26238 34130
rect 26290 34078 26292 34130
rect 26236 34066 26292 34078
rect 26348 33908 26404 33918
rect 26348 33234 26404 33852
rect 26572 33796 26628 34862
rect 27020 34802 27076 35868
rect 27132 35588 27188 35598
rect 27132 35364 27188 35532
rect 27132 35298 27188 35308
rect 27132 35028 27188 35038
rect 27132 34914 27188 34972
rect 27132 34862 27134 34914
rect 27186 34862 27188 34914
rect 27132 34850 27188 34862
rect 27020 34750 27022 34802
rect 27074 34750 27076 34802
rect 27020 34692 27076 34750
rect 27020 34626 27076 34636
rect 27244 34468 27300 36988
rect 27020 34412 27300 34468
rect 27356 37940 27412 37950
rect 27356 37042 27412 37884
rect 27580 37828 27636 38612
rect 28140 38612 28196 38668
rect 28252 38724 28308 38734
rect 28476 38722 28532 39564
rect 28476 38670 28478 38722
rect 28530 38670 28532 38722
rect 28252 38612 28420 38668
rect 28140 38546 28196 38556
rect 28028 38500 28084 38510
rect 27356 36990 27358 37042
rect 27410 36990 27412 37042
rect 27020 34132 27076 34412
rect 27020 34076 27188 34132
rect 26348 33182 26350 33234
rect 26402 33182 26404 33234
rect 26348 33170 26404 33182
rect 26460 33684 26516 33694
rect 26012 32676 26068 32686
rect 25788 31218 25956 31220
rect 25788 31166 25790 31218
rect 25842 31166 25956 31218
rect 25788 31164 25956 31166
rect 25788 31154 25844 31164
rect 25900 30660 25956 31164
rect 26012 30994 26068 32620
rect 26348 32564 26404 32574
rect 26460 32564 26516 33628
rect 26348 32562 26516 32564
rect 26348 32510 26350 32562
rect 26402 32510 26516 32562
rect 26348 32508 26516 32510
rect 26348 32498 26404 32508
rect 26012 30942 26014 30994
rect 26066 30942 26068 30994
rect 26012 30930 26068 30942
rect 26460 31220 26516 31230
rect 26572 31220 26628 33740
rect 26796 33572 26852 33582
rect 26796 33478 26852 33516
rect 27020 33348 27076 33358
rect 26908 33236 26964 33246
rect 26796 32338 26852 32350
rect 26796 32286 26798 32338
rect 26850 32286 26852 32338
rect 26796 31778 26852 32286
rect 26796 31726 26798 31778
rect 26850 31726 26852 31778
rect 26460 31218 26628 31220
rect 26460 31166 26462 31218
rect 26514 31166 26628 31218
rect 26460 31164 26628 31166
rect 26684 31444 26740 31454
rect 26684 31218 26740 31388
rect 26684 31166 26686 31218
rect 26738 31166 26740 31218
rect 26348 30884 26404 30894
rect 25900 30604 26180 30660
rect 26012 30436 26068 30446
rect 25676 30434 26068 30436
rect 25676 30382 26014 30434
rect 26066 30382 26068 30434
rect 25676 30380 26068 30382
rect 26012 30370 26068 30380
rect 25452 30210 25508 30222
rect 25788 30212 25844 30222
rect 26124 30212 26180 30604
rect 25452 30158 25454 30210
rect 25506 30158 25508 30210
rect 25452 30100 25508 30158
rect 25452 30034 25508 30044
rect 25564 30156 25788 30212
rect 25564 29650 25620 30156
rect 25788 30146 25844 30156
rect 26012 30156 26180 30212
rect 26348 30210 26404 30828
rect 26348 30158 26350 30210
rect 26402 30158 26404 30210
rect 25900 30100 25956 30110
rect 25900 30006 25956 30044
rect 26012 29652 26068 30156
rect 26348 30146 26404 30158
rect 26460 30212 26516 31164
rect 26684 31154 26740 31166
rect 26796 30996 26852 31726
rect 26796 30930 26852 30940
rect 26460 30146 26516 30156
rect 26572 30882 26628 30894
rect 26572 30830 26574 30882
rect 26626 30830 26628 30882
rect 26572 30210 26628 30830
rect 26572 30158 26574 30210
rect 26626 30158 26628 30210
rect 26572 30146 26628 30158
rect 26908 30100 26964 33180
rect 27020 31668 27076 33292
rect 27132 31890 27188 34076
rect 27244 34020 27300 34030
rect 27244 33684 27300 33964
rect 27244 33618 27300 33628
rect 27244 33236 27300 33246
rect 27356 33236 27412 36990
rect 27468 37604 27524 37614
rect 27468 35810 27524 37548
rect 27580 37266 27636 37772
rect 27580 37214 27582 37266
rect 27634 37214 27636 37266
rect 27580 37202 27636 37214
rect 27916 38388 27972 38398
rect 27804 37156 27860 37166
rect 27804 37062 27860 37100
rect 27580 36596 27636 36606
rect 27580 36502 27636 36540
rect 27916 36372 27972 38332
rect 28028 37490 28084 38444
rect 28364 38162 28420 38612
rect 28364 38110 28366 38162
rect 28418 38110 28420 38162
rect 28364 38098 28420 38110
rect 28252 38050 28308 38062
rect 28252 37998 28254 38050
rect 28306 37998 28308 38050
rect 28140 37940 28196 37950
rect 28252 37940 28308 37998
rect 28476 37940 28532 38670
rect 28588 38276 28644 39788
rect 28700 39842 28756 40124
rect 28700 39790 28702 39842
rect 28754 39790 28756 39842
rect 28700 39778 28756 39790
rect 29036 38724 29092 38734
rect 29036 38630 29092 38668
rect 29372 38668 29428 40796
rect 29820 40292 29876 40302
rect 29820 40198 29876 40236
rect 29596 40068 29652 40078
rect 29596 39730 29652 40012
rect 29596 39678 29598 39730
rect 29650 39678 29652 39730
rect 29596 39666 29652 39678
rect 29932 39620 29988 42140
rect 30156 41972 30212 41982
rect 30268 41972 30324 43484
rect 30716 43316 30772 43326
rect 30156 41970 30324 41972
rect 30156 41918 30158 41970
rect 30210 41918 30324 41970
rect 30156 41916 30324 41918
rect 30156 41906 30212 41916
rect 30156 41524 30212 41534
rect 30156 41298 30212 41468
rect 30156 41246 30158 41298
rect 30210 41246 30212 41298
rect 30156 41234 30212 41246
rect 30268 40068 30324 41916
rect 30380 43314 30772 43316
rect 30380 43262 30718 43314
rect 30770 43262 30772 43314
rect 30380 43260 30772 43262
rect 30380 42866 30436 43260
rect 30716 43250 30772 43260
rect 30380 42814 30382 42866
rect 30434 42814 30436 42866
rect 30380 41410 30436 42814
rect 30604 42756 30660 42766
rect 30492 42420 30548 42430
rect 30492 41860 30548 42364
rect 30604 42082 30660 42700
rect 30716 42756 30772 42766
rect 30828 42756 30884 44270
rect 30940 43650 30996 43662
rect 30940 43598 30942 43650
rect 30994 43598 30996 43650
rect 30940 43540 30996 43598
rect 30940 43474 30996 43484
rect 30716 42754 30884 42756
rect 30716 42702 30718 42754
rect 30770 42702 30884 42754
rect 30716 42700 30884 42702
rect 31052 43314 31108 43326
rect 31052 43262 31054 43314
rect 31106 43262 31108 43314
rect 31052 42756 31108 43262
rect 31164 42756 31220 42766
rect 31052 42754 31220 42756
rect 31052 42702 31166 42754
rect 31218 42702 31220 42754
rect 31052 42700 31220 42702
rect 30716 42690 30772 42700
rect 31164 42690 31220 42700
rect 30604 42030 30606 42082
rect 30658 42030 30660 42082
rect 30604 42018 30660 42030
rect 30940 42642 30996 42654
rect 30940 42590 30942 42642
rect 30994 42590 30996 42642
rect 30940 41860 30996 42590
rect 30492 41804 30660 41860
rect 30380 41358 30382 41410
rect 30434 41358 30436 41410
rect 30380 41346 30436 41358
rect 30492 41186 30548 41198
rect 30492 41134 30494 41186
rect 30546 41134 30548 41186
rect 30492 40404 30548 41134
rect 30492 40310 30548 40348
rect 30268 40012 30436 40068
rect 30268 39844 30324 39854
rect 30268 39750 30324 39788
rect 30156 39620 30212 39630
rect 30380 39620 30436 40012
rect 29708 39618 30212 39620
rect 29708 39566 30158 39618
rect 30210 39566 30212 39618
rect 29708 39564 30212 39566
rect 29596 39060 29652 39070
rect 29708 39060 29764 39564
rect 30156 39554 30212 39564
rect 30268 39564 30436 39620
rect 29596 39058 29764 39060
rect 29596 39006 29598 39058
rect 29650 39006 29764 39058
rect 29596 39004 29764 39006
rect 29596 38994 29652 39004
rect 29372 38612 29988 38668
rect 28588 38210 28644 38220
rect 29260 38388 29316 38398
rect 29260 38162 29316 38332
rect 29260 38110 29262 38162
rect 29314 38110 29316 38162
rect 29260 38098 29316 38110
rect 28196 37884 28308 37940
rect 28364 37884 28532 37940
rect 28588 38050 28644 38062
rect 28588 37998 28590 38050
rect 28642 37998 28644 38050
rect 28140 37874 28196 37884
rect 28364 37604 28420 37884
rect 28028 37438 28030 37490
rect 28082 37438 28084 37490
rect 28028 37426 28084 37438
rect 28140 37548 28420 37604
rect 28476 37604 28532 37614
rect 28028 36372 28084 36382
rect 27916 36316 28028 36372
rect 28028 36258 28084 36316
rect 28028 36206 28030 36258
rect 28082 36206 28084 36258
rect 27468 35758 27470 35810
rect 27522 35758 27524 35810
rect 27468 33684 27524 35758
rect 27580 35812 27636 35822
rect 27580 34914 27636 35756
rect 27804 35700 27860 35710
rect 27804 35606 27860 35644
rect 27580 34862 27582 34914
rect 27634 34862 27636 34914
rect 27580 34132 27636 34862
rect 27804 35364 27860 35374
rect 27804 34914 27860 35308
rect 28028 35364 28084 36206
rect 28028 35298 28084 35308
rect 28140 35140 28196 37548
rect 28476 37492 28532 37548
rect 28252 37436 28532 37492
rect 28252 37378 28308 37436
rect 28252 37326 28254 37378
rect 28306 37326 28308 37378
rect 28252 37314 28308 37326
rect 28364 37266 28420 37278
rect 28364 37214 28366 37266
rect 28418 37214 28420 37266
rect 28364 36372 28420 37214
rect 28476 37156 28532 37166
rect 28588 37156 28644 37998
rect 29820 38050 29876 38062
rect 29820 37998 29822 38050
rect 29874 37998 29876 38050
rect 28532 37100 28644 37156
rect 28700 37940 28756 37950
rect 28476 37090 28532 37100
rect 28700 36482 28756 37884
rect 29708 37828 29764 37838
rect 29708 37734 29764 37772
rect 29036 37492 29092 37502
rect 29036 37398 29092 37436
rect 29484 37492 29540 37502
rect 29484 37398 29540 37436
rect 29708 37492 29764 37502
rect 29820 37492 29876 37998
rect 29708 37490 29876 37492
rect 29708 37438 29710 37490
rect 29762 37438 29876 37490
rect 29708 37436 29876 37438
rect 29708 37426 29764 37436
rect 29596 37380 29652 37390
rect 29596 37286 29652 37324
rect 28700 36430 28702 36482
rect 28754 36430 28756 36482
rect 28700 36418 28756 36430
rect 28924 37268 28980 37278
rect 28364 36278 28420 36316
rect 28476 36260 28532 36270
rect 28476 36166 28532 36204
rect 28700 35924 28756 35934
rect 28700 35830 28756 35868
rect 28252 35700 28308 35710
rect 28252 35606 28308 35644
rect 28140 35074 28196 35084
rect 27804 34862 27806 34914
rect 27858 34862 27860 34914
rect 27804 34850 27860 34862
rect 28252 34916 28308 34926
rect 28308 34860 28420 34916
rect 28252 34822 28308 34860
rect 27692 34692 27748 34702
rect 27692 34598 27748 34636
rect 28140 34692 28196 34702
rect 28364 34692 28420 34860
rect 28700 34692 28756 34702
rect 28364 34690 28756 34692
rect 28364 34638 28702 34690
rect 28754 34638 28756 34690
rect 28364 34636 28756 34638
rect 28924 34692 28980 37212
rect 29820 37268 29876 37278
rect 29820 37174 29876 37212
rect 29596 37156 29652 37166
rect 29148 36708 29204 36718
rect 29148 35922 29204 36652
rect 29260 36260 29316 36270
rect 29260 36166 29316 36204
rect 29148 35870 29150 35922
rect 29202 35870 29204 35922
rect 29148 35364 29204 35870
rect 29148 35298 29204 35308
rect 29036 35140 29092 35150
rect 29036 34914 29092 35084
rect 29036 34862 29038 34914
rect 29090 34862 29092 34914
rect 29036 34850 29092 34862
rect 29372 34802 29428 34814
rect 29372 34750 29374 34802
rect 29426 34750 29428 34802
rect 29260 34692 29316 34702
rect 28924 34636 29092 34692
rect 28028 34244 28084 34254
rect 27916 34188 28028 34244
rect 27580 34076 27748 34132
rect 27580 33908 27636 33918
rect 27580 33814 27636 33852
rect 27468 33628 27636 33684
rect 27300 33180 27412 33236
rect 27244 33170 27300 33180
rect 27468 32900 27524 32910
rect 27468 32562 27524 32844
rect 27580 32676 27636 33628
rect 27692 33572 27748 34076
rect 27692 33506 27748 33516
rect 27804 34020 27860 34030
rect 27804 33346 27860 33964
rect 27916 33458 27972 34188
rect 28028 34150 28084 34188
rect 28140 34242 28196 34636
rect 28140 34190 28142 34242
rect 28194 34190 28196 34242
rect 28140 34178 28196 34190
rect 28252 34580 28308 34590
rect 28252 34242 28308 34524
rect 28252 34190 28254 34242
rect 28306 34190 28308 34242
rect 28252 34020 28308 34190
rect 28252 33954 28308 33964
rect 28700 33908 28756 34636
rect 28700 33842 28756 33852
rect 28812 34018 28868 34030
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 27916 33406 27918 33458
rect 27970 33406 27972 33458
rect 27916 33394 27972 33406
rect 28476 33572 28532 33582
rect 27804 33294 27806 33346
rect 27858 33294 27860 33346
rect 27804 33282 27860 33294
rect 28028 33348 28084 33358
rect 28028 33254 28084 33292
rect 28252 33236 28308 33246
rect 28252 33142 28308 33180
rect 27580 32610 27636 32620
rect 27692 33124 27748 33134
rect 27468 32510 27470 32562
rect 27522 32510 27524 32562
rect 27468 32498 27524 32510
rect 27692 32340 27748 33068
rect 28476 32788 28532 33516
rect 28812 33348 28868 33966
rect 28812 33282 28868 33292
rect 28924 32788 28980 32798
rect 28476 32786 28980 32788
rect 28476 32734 28926 32786
rect 28978 32734 28980 32786
rect 28476 32732 28980 32734
rect 28364 32676 28420 32686
rect 28364 32582 28420 32620
rect 28476 32674 28532 32732
rect 28924 32722 28980 32732
rect 28476 32622 28478 32674
rect 28530 32622 28532 32674
rect 28476 32610 28532 32622
rect 28140 32564 28196 32574
rect 27692 32274 27748 32284
rect 27804 32562 28196 32564
rect 27804 32510 28142 32562
rect 28194 32510 28196 32562
rect 27804 32508 28196 32510
rect 27132 31838 27134 31890
rect 27186 31838 27188 31890
rect 27132 31826 27188 31838
rect 27356 31780 27412 31790
rect 27356 31778 27748 31780
rect 27356 31726 27358 31778
rect 27410 31726 27748 31778
rect 27356 31724 27748 31726
rect 27356 31714 27412 31724
rect 27020 31612 27300 31668
rect 27020 30322 27076 31612
rect 27020 30270 27022 30322
rect 27074 30270 27076 30322
rect 27020 30258 27076 30270
rect 27132 31332 27188 31342
rect 26908 30044 27076 30100
rect 25564 29598 25566 29650
rect 25618 29598 25620 29650
rect 25564 29586 25620 29598
rect 25900 29650 26068 29652
rect 25900 29598 26014 29650
rect 26066 29598 26068 29650
rect 25900 29596 26068 29598
rect 25788 29202 25844 29214
rect 25788 29150 25790 29202
rect 25842 29150 25844 29202
rect 25452 28420 25508 28430
rect 25452 28084 25508 28364
rect 25452 28082 25620 28084
rect 25452 28030 25454 28082
rect 25506 28030 25620 28082
rect 25452 28028 25620 28030
rect 25452 28018 25508 28028
rect 25564 26964 25620 28028
rect 25788 28082 25844 29150
rect 25900 28420 25956 29596
rect 26012 29586 26068 29596
rect 26124 29986 26180 29998
rect 26124 29934 26126 29986
rect 26178 29934 26180 29986
rect 26124 29202 26180 29934
rect 26124 29150 26126 29202
rect 26178 29150 26180 29202
rect 26124 29138 26180 29150
rect 26684 29314 26740 29326
rect 26684 29262 26686 29314
rect 26738 29262 26740 29314
rect 26348 29092 26404 29102
rect 26236 28980 26292 28990
rect 26012 28924 26236 28980
rect 26012 28644 26068 28924
rect 26236 28914 26292 28924
rect 26348 28756 26404 29036
rect 26684 28868 26740 29262
rect 26684 28802 26740 28812
rect 26908 28980 26964 28990
rect 26348 28754 26516 28756
rect 26348 28702 26350 28754
rect 26402 28702 26516 28754
rect 26348 28700 26516 28702
rect 26348 28690 26404 28700
rect 26012 28550 26068 28588
rect 25900 28364 26068 28420
rect 25788 28030 25790 28082
rect 25842 28030 25844 28082
rect 25788 28018 25844 28030
rect 25676 27858 25732 27870
rect 25676 27806 25678 27858
rect 25730 27806 25732 27858
rect 25676 27748 25732 27806
rect 25676 27682 25732 27692
rect 25900 27858 25956 27870
rect 25900 27806 25902 27858
rect 25954 27806 25956 27858
rect 25900 27636 25956 27806
rect 25900 27076 25956 27580
rect 25900 27010 25956 27020
rect 26012 27074 26068 28364
rect 26460 27860 26516 28700
rect 26908 28754 26964 28924
rect 26908 28702 26910 28754
rect 26962 28702 26964 28754
rect 26908 28690 26964 28702
rect 27020 28082 27076 30044
rect 27020 28030 27022 28082
rect 27074 28030 27076 28082
rect 27020 28018 27076 28030
rect 26460 27766 26516 27804
rect 26684 27972 26740 27982
rect 26684 27636 26740 27916
rect 27132 27860 27188 31276
rect 27244 30994 27300 31612
rect 27692 31220 27748 31724
rect 27804 31666 27860 32508
rect 28140 32498 28196 32508
rect 27804 31614 27806 31666
rect 27858 31614 27860 31666
rect 27804 31602 27860 31614
rect 28028 31668 28084 31678
rect 28028 31574 28084 31612
rect 28476 31444 28532 31454
rect 27804 31220 27860 31230
rect 27692 31218 27860 31220
rect 27692 31166 27806 31218
rect 27858 31166 27860 31218
rect 27692 31164 27860 31166
rect 27804 31154 27860 31164
rect 28476 31220 28532 31388
rect 28812 31220 28868 31230
rect 28476 31218 28868 31220
rect 28476 31166 28478 31218
rect 28530 31166 28814 31218
rect 28866 31166 28868 31218
rect 28476 31164 28868 31166
rect 28476 31154 28532 31164
rect 28812 31154 28868 31164
rect 29036 31218 29092 34636
rect 29260 34598 29316 34636
rect 29372 34244 29428 34750
rect 29372 34178 29428 34188
rect 29260 34020 29316 34030
rect 29260 33926 29316 33964
rect 29484 34020 29540 34030
rect 29260 33236 29316 33246
rect 29148 33124 29204 33134
rect 29148 31890 29204 33068
rect 29148 31838 29150 31890
rect 29202 31838 29204 31890
rect 29148 31826 29204 31838
rect 29036 31166 29038 31218
rect 29090 31166 29092 31218
rect 29036 31154 29092 31166
rect 27244 30942 27246 30994
rect 27298 30942 27300 30994
rect 27244 30930 27300 30942
rect 27692 30996 27748 31006
rect 27692 30902 27748 30940
rect 27916 30994 27972 31006
rect 27916 30942 27918 30994
rect 27970 30942 27972 30994
rect 27916 30772 27972 30942
rect 27916 30548 27972 30716
rect 28924 30882 28980 30894
rect 28924 30830 28926 30882
rect 28978 30830 28980 30882
rect 27916 30492 28196 30548
rect 28028 30212 28084 30222
rect 27244 29652 27300 29662
rect 27244 29558 27300 29596
rect 27804 29652 27860 29662
rect 27804 29558 27860 29596
rect 27468 29540 27524 29550
rect 27468 28754 27524 29484
rect 27580 29538 27636 29550
rect 27580 29486 27582 29538
rect 27634 29486 27636 29538
rect 27580 28868 27636 29486
rect 27916 29540 27972 29550
rect 27916 29446 27972 29484
rect 27580 28802 27636 28812
rect 28028 29426 28084 30156
rect 28140 30100 28196 30492
rect 28588 30212 28644 30222
rect 28588 30118 28644 30156
rect 28140 30006 28196 30044
rect 28924 29652 28980 30830
rect 28924 29596 29092 29652
rect 28588 29540 28644 29550
rect 28644 29484 28756 29540
rect 28588 29446 28644 29484
rect 28028 29374 28030 29426
rect 28082 29374 28084 29426
rect 28028 28756 28084 29374
rect 28364 29428 28420 29438
rect 28364 29334 28420 29372
rect 28700 29092 28756 29484
rect 28700 29026 28756 29036
rect 28924 29426 28980 29438
rect 28924 29374 28926 29426
rect 28978 29374 28980 29426
rect 28812 28868 28868 28878
rect 28924 28868 28980 29374
rect 29036 29428 29092 29596
rect 29260 29540 29316 33180
rect 29484 30996 29540 33964
rect 29596 33796 29652 37100
rect 29708 36484 29764 36494
rect 29708 36390 29764 36428
rect 29820 34804 29876 34814
rect 29820 34710 29876 34748
rect 29932 34468 29988 38612
rect 30044 38164 30100 38174
rect 30044 38070 30100 38108
rect 30044 37266 30100 37278
rect 30044 37214 30046 37266
rect 30098 37214 30100 37266
rect 30044 37156 30100 37214
rect 30044 37090 30100 37100
rect 30156 35924 30212 35934
rect 30044 35868 30156 35924
rect 30044 34804 30100 35868
rect 30156 35858 30212 35868
rect 30044 34738 30100 34748
rect 30156 34692 30212 34702
rect 30156 34598 30212 34636
rect 29820 34412 29988 34468
rect 29820 34244 29876 34412
rect 29820 34188 30212 34244
rect 29932 34020 29988 34030
rect 29932 33926 29988 33964
rect 29596 33740 29988 33796
rect 29708 31556 29764 31566
rect 29708 31220 29764 31500
rect 29708 31154 29764 31164
rect 29484 30902 29540 30940
rect 29260 29484 29428 29540
rect 29036 29362 29092 29372
rect 28868 28812 28980 28868
rect 28812 28802 28868 28812
rect 27468 28702 27470 28754
rect 27522 28702 27524 28754
rect 27468 28644 27524 28702
rect 27468 28578 27524 28588
rect 27916 28700 28084 28756
rect 29260 28756 29316 28766
rect 27580 28532 27636 28542
rect 27356 27972 27412 27982
rect 27356 27878 27412 27916
rect 26684 27542 26740 27580
rect 27020 27804 27188 27860
rect 27580 27858 27636 28476
rect 27580 27806 27582 27858
rect 27634 27806 27636 27858
rect 26012 27022 26014 27074
rect 26066 27022 26068 27074
rect 25788 26964 25844 26974
rect 25564 26962 25844 26964
rect 25564 26910 25790 26962
rect 25842 26910 25844 26962
rect 25564 26908 25844 26910
rect 25788 26898 25844 26908
rect 26012 26516 26068 27022
rect 26572 26850 26628 26862
rect 26572 26798 26574 26850
rect 26626 26798 26628 26850
rect 26572 26516 26628 26798
rect 27020 26628 27076 27804
rect 27132 27188 27188 27198
rect 27580 27188 27636 27806
rect 27132 27186 27636 27188
rect 27132 27134 27134 27186
rect 27186 27134 27636 27186
rect 27132 27132 27636 27134
rect 27132 27122 27188 27132
rect 27916 26908 27972 28700
rect 28364 28644 28420 28654
rect 28252 28530 28308 28542
rect 28252 28478 28254 28530
rect 28306 28478 28308 28530
rect 27020 26562 27076 26572
rect 27804 26852 27972 26908
rect 28028 28420 28084 28430
rect 28252 28420 28308 28478
rect 28364 28530 28420 28588
rect 28588 28644 28644 28654
rect 28588 28550 28644 28588
rect 29148 28644 29204 28654
rect 29148 28550 29204 28588
rect 29260 28642 29316 28700
rect 29260 28590 29262 28642
rect 29314 28590 29316 28642
rect 29260 28578 29316 28590
rect 28364 28478 28366 28530
rect 28418 28478 28420 28530
rect 28364 28466 28420 28478
rect 28028 28418 28308 28420
rect 28028 28366 28030 28418
rect 28082 28366 28308 28418
rect 28028 28364 28308 28366
rect 26012 26514 26628 26516
rect 26012 26462 26014 26514
rect 26066 26462 26574 26514
rect 26626 26462 26628 26514
rect 26012 26460 26628 26462
rect 26012 26450 26068 26460
rect 26572 26450 26628 26460
rect 27804 26404 27860 26852
rect 25396 26348 25620 26404
rect 25340 26310 25396 26348
rect 25228 26180 25284 26236
rect 25452 26180 25508 26190
rect 25228 26178 25508 26180
rect 25228 26126 25454 26178
rect 25506 26126 25508 26178
rect 25228 26124 25508 26126
rect 25452 26114 25508 26124
rect 25228 25956 25284 25966
rect 25228 25620 25284 25900
rect 25228 25506 25284 25564
rect 25228 25454 25230 25506
rect 25282 25454 25284 25506
rect 25228 25442 25284 25454
rect 25564 25506 25620 26348
rect 27804 26338 27860 26348
rect 27132 25620 27188 25630
rect 27132 25526 27188 25564
rect 25564 25454 25566 25506
rect 25618 25454 25620 25506
rect 25564 25442 25620 25454
rect 27916 25508 27972 25518
rect 25004 24836 25060 24846
rect 25060 24780 25172 24836
rect 25004 24770 25060 24780
rect 25116 24052 25172 24780
rect 25788 24722 25844 24734
rect 25788 24670 25790 24722
rect 25842 24670 25844 24722
rect 25340 24610 25396 24622
rect 25788 24612 25844 24670
rect 25340 24558 25342 24610
rect 25394 24558 25396 24610
rect 25228 24052 25284 24062
rect 25116 24050 25284 24052
rect 25116 23998 25230 24050
rect 25282 23998 25284 24050
rect 25116 23996 25284 23998
rect 25228 23986 25284 23996
rect 24780 23940 24836 23950
rect 24780 23846 24836 23884
rect 24556 23762 24612 23772
rect 25228 23828 25284 23838
rect 25340 23828 25396 24558
rect 25284 23772 25396 23828
rect 25452 24556 25788 24612
rect 25452 23940 25508 24556
rect 25788 24546 25844 24556
rect 26236 24612 26292 24622
rect 26236 24518 26292 24556
rect 27916 24276 27972 25452
rect 27916 24210 27972 24220
rect 25788 24052 25844 24062
rect 25788 23958 25844 23996
rect 25228 23762 25284 23772
rect 22988 23378 23156 23380
rect 22988 23326 22990 23378
rect 23042 23326 23156 23378
rect 22988 23324 23156 23326
rect 25452 23378 25508 23884
rect 25452 23326 25454 23378
rect 25506 23326 25508 23378
rect 22204 23268 22260 23278
rect 21980 23212 22204 23268
rect 21308 23174 21364 23212
rect 22204 23174 22260 23212
rect 22988 23268 23044 23324
rect 25452 23314 25508 23326
rect 22988 23202 23044 23212
rect 19068 22930 19348 22932
rect 19068 22878 19070 22930
rect 19122 22878 19348 22930
rect 19068 22876 19348 22878
rect 28028 22932 28084 28364
rect 28252 27972 28308 28364
rect 28252 27906 28308 27916
rect 28140 27860 28196 27870
rect 28140 27766 28196 27804
rect 29372 27858 29428 29484
rect 29596 29426 29652 29438
rect 29596 29374 29598 29426
rect 29650 29374 29652 29426
rect 29484 29092 29540 29102
rect 29484 28642 29540 29036
rect 29484 28590 29486 28642
rect 29538 28590 29540 28642
rect 29484 28578 29540 28590
rect 29596 28644 29652 29374
rect 29596 28578 29652 28588
rect 29708 29428 29764 29438
rect 29708 28642 29764 29372
rect 29932 29202 29988 33740
rect 29932 29150 29934 29202
rect 29986 29150 29988 29202
rect 29932 29138 29988 29150
rect 30156 28866 30212 34188
rect 30268 33572 30324 39564
rect 30380 39396 30436 39406
rect 30380 34916 30436 39340
rect 30604 38836 30660 41804
rect 30940 41794 30996 41804
rect 31388 41188 31444 41198
rect 31388 41094 31444 41132
rect 31164 41076 31220 41086
rect 31164 40982 31220 41020
rect 30828 40402 30884 40414
rect 30828 40350 30830 40402
rect 30882 40350 30884 40402
rect 30828 40068 30884 40350
rect 31164 40402 31220 40414
rect 31164 40350 31166 40402
rect 31218 40350 31220 40402
rect 30884 40012 30996 40068
rect 30828 40002 30884 40012
rect 30716 39618 30772 39630
rect 30716 39566 30718 39618
rect 30770 39566 30772 39618
rect 30716 38948 30772 39566
rect 30940 39618 30996 40012
rect 30940 39566 30942 39618
rect 30994 39566 30996 39618
rect 30940 39554 30996 39566
rect 30940 38948 30996 38958
rect 30716 38946 30996 38948
rect 30716 38894 30942 38946
rect 30994 38894 30996 38946
rect 30716 38892 30996 38894
rect 30940 38882 30996 38892
rect 30604 38780 30884 38836
rect 30828 38668 30884 38780
rect 30492 38612 30548 38622
rect 30492 38050 30548 38556
rect 30492 37998 30494 38050
rect 30546 37998 30548 38050
rect 30492 37986 30548 37998
rect 30716 38612 30884 38668
rect 31164 38724 31220 40350
rect 31612 39844 31668 47068
rect 31724 43652 31780 48076
rect 32172 48130 32228 48188
rect 32172 48078 32174 48130
rect 32226 48078 32228 48130
rect 32060 47572 32116 47582
rect 32060 47478 32116 47516
rect 31948 46788 32004 46798
rect 31836 45892 31892 45902
rect 31836 45798 31892 45836
rect 31724 43558 31780 43596
rect 31612 39788 31780 39844
rect 31388 39618 31444 39630
rect 31388 39566 31390 39618
rect 31442 39566 31444 39618
rect 31388 38948 31444 39566
rect 31724 39060 31780 39788
rect 31724 38994 31780 39004
rect 31836 39618 31892 39630
rect 31836 39566 31838 39618
rect 31890 39566 31892 39618
rect 31388 38892 31556 38948
rect 31276 38836 31332 38846
rect 31276 38834 31444 38836
rect 31276 38782 31278 38834
rect 31330 38782 31444 38834
rect 31276 38780 31444 38782
rect 31276 38770 31332 38780
rect 31164 38658 31220 38668
rect 31052 38612 31108 38622
rect 30604 37940 30660 37950
rect 30604 37846 30660 37884
rect 30492 37044 30548 37054
rect 30492 36950 30548 36988
rect 30380 34850 30436 34860
rect 30604 35364 30660 35374
rect 30380 34692 30436 34702
rect 30380 34130 30436 34636
rect 30380 34078 30382 34130
rect 30434 34078 30436 34130
rect 30380 34066 30436 34078
rect 30268 33506 30324 33516
rect 30492 33908 30548 33918
rect 30380 33346 30436 33358
rect 30380 33294 30382 33346
rect 30434 33294 30436 33346
rect 30380 29652 30436 33294
rect 30492 31890 30548 33852
rect 30492 31838 30494 31890
rect 30546 31838 30548 31890
rect 30492 31826 30548 31838
rect 30380 29586 30436 29596
rect 30492 30324 30548 30334
rect 30604 30324 30660 35308
rect 30492 30322 30660 30324
rect 30492 30270 30494 30322
rect 30546 30270 30660 30322
rect 30492 30268 30660 30270
rect 30492 28980 30548 30268
rect 30716 29988 30772 38612
rect 31052 37266 31108 38556
rect 31388 38500 31444 38780
rect 31388 38434 31444 38444
rect 31052 37214 31054 37266
rect 31106 37214 31108 37266
rect 31052 37202 31108 37214
rect 31164 38388 31220 38398
rect 30828 35252 30884 35262
rect 30828 34130 30884 35196
rect 31052 34916 31108 34926
rect 30940 34692 30996 34702
rect 30940 34598 30996 34636
rect 30828 34078 30830 34130
rect 30882 34078 30884 34130
rect 30828 34066 30884 34078
rect 30940 33124 30996 33134
rect 30940 33030 30996 33068
rect 30940 31556 30996 31566
rect 30940 30212 30996 31500
rect 30940 30118 30996 30156
rect 30716 29922 30772 29932
rect 30492 28914 30548 28924
rect 30156 28814 30158 28866
rect 30210 28814 30212 28866
rect 30156 28802 30212 28814
rect 29708 28590 29710 28642
rect 29762 28590 29764 28642
rect 29708 28578 29764 28590
rect 31052 28308 31108 34860
rect 31052 28242 31108 28252
rect 31164 28196 31220 38332
rect 31276 38164 31332 38174
rect 31276 37266 31332 38108
rect 31500 37604 31556 38892
rect 31724 38834 31780 38846
rect 31724 38782 31726 38834
rect 31778 38782 31780 38834
rect 31724 37828 31780 38782
rect 31836 38050 31892 39566
rect 31948 38836 32004 46732
rect 32060 46004 32116 46014
rect 32060 45910 32116 45948
rect 32172 45332 32228 48078
rect 32172 45266 32228 45276
rect 32508 47012 32564 47022
rect 32508 45108 32564 46956
rect 32620 46898 32676 51212
rect 33180 52162 33572 52164
rect 33180 52110 33406 52162
rect 33458 52110 33572 52162
rect 33180 52108 33572 52110
rect 33180 50036 33236 52108
rect 33404 52098 33460 52108
rect 34636 50708 34692 53564
rect 34748 52164 34804 54350
rect 36092 54404 36148 54414
rect 36092 54310 36148 54348
rect 36428 54290 36484 55358
rect 37100 55298 37156 56142
rect 39788 56194 39844 56206
rect 39788 56142 39790 56194
rect 39842 56142 39844 56194
rect 38892 55970 38948 55982
rect 38892 55918 38894 55970
rect 38946 55918 38948 55970
rect 38892 55860 38948 55918
rect 38892 55794 38948 55804
rect 39788 55468 39844 56142
rect 40124 56194 40180 56590
rect 41020 56308 41076 59200
rect 41468 56308 41524 56318
rect 41020 56306 41524 56308
rect 41020 56254 41470 56306
rect 41522 56254 41524 56306
rect 41020 56252 41524 56254
rect 41468 56242 41524 56252
rect 43260 56308 43316 59200
rect 43260 56242 43316 56252
rect 44604 56308 44660 56318
rect 44604 56214 44660 56252
rect 40124 56142 40126 56194
rect 40178 56142 40180 56194
rect 40124 56130 40180 56142
rect 40460 56082 40516 56094
rect 40460 56030 40462 56082
rect 40514 56030 40516 56082
rect 40460 55860 40516 56030
rect 40460 55794 40516 55804
rect 43708 56082 43764 56094
rect 43708 56030 43710 56082
rect 43762 56030 43764 56082
rect 39116 55412 39844 55468
rect 43148 55412 43204 55422
rect 39116 55410 39172 55412
rect 39116 55358 39118 55410
rect 39170 55358 39172 55410
rect 39116 55346 39172 55358
rect 42924 55410 43204 55412
rect 42924 55358 43150 55410
rect 43202 55358 43204 55410
rect 42924 55356 43204 55358
rect 37100 55246 37102 55298
rect 37154 55246 37156 55298
rect 37100 55234 37156 55246
rect 38332 55298 38388 55310
rect 38332 55246 38334 55298
rect 38386 55246 38388 55298
rect 37324 55186 37380 55198
rect 37324 55134 37326 55186
rect 37378 55134 37380 55186
rect 36428 54238 36430 54290
rect 36482 54238 36484 54290
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 36428 53058 36484 54238
rect 36876 54628 36932 54638
rect 36876 54402 36932 54572
rect 36876 54350 36878 54402
rect 36930 54350 36932 54402
rect 36764 53732 36820 53742
rect 36428 53006 36430 53058
rect 36482 53006 36484 53058
rect 36428 52994 36484 53006
rect 36540 53060 36596 53070
rect 36540 52966 36596 53004
rect 36764 52946 36820 53676
rect 36764 52894 36766 52946
rect 36818 52894 36820 52946
rect 36764 52882 36820 52894
rect 35980 52836 36036 52846
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34860 52164 34916 52174
rect 34748 52108 34860 52164
rect 34860 52098 34916 52108
rect 35980 52164 36036 52780
rect 36204 52834 36260 52846
rect 36204 52782 36206 52834
rect 36258 52782 36260 52834
rect 36204 52276 36260 52782
rect 36204 52182 36260 52220
rect 36316 52500 36372 52510
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 34636 50706 35252 50708
rect 34636 50654 34638 50706
rect 34690 50654 35252 50706
rect 34636 50652 35252 50654
rect 34636 50642 34692 50652
rect 35196 50594 35252 50652
rect 35196 50542 35198 50594
rect 35250 50542 35252 50594
rect 35196 50530 35252 50542
rect 33180 49942 33236 49980
rect 34972 50370 35028 50382
rect 34972 50318 34974 50370
rect 35026 50318 35028 50370
rect 34412 49698 34468 49710
rect 34412 49646 34414 49698
rect 34466 49646 34468 49698
rect 32844 49252 32900 49262
rect 32844 49028 32900 49196
rect 34188 49252 34244 49262
rect 32620 46846 32622 46898
rect 32674 46846 32676 46898
rect 32620 46452 32676 46846
rect 32620 46386 32676 46396
rect 32732 49026 32900 49028
rect 32732 48974 32846 49026
rect 32898 48974 32900 49026
rect 32732 48972 32900 48974
rect 32732 45890 32788 48972
rect 32844 48962 32900 48972
rect 33068 49140 33124 49150
rect 33068 48914 33124 49084
rect 34188 49026 34244 49196
rect 34188 48974 34190 49026
rect 34242 48974 34244 49026
rect 34188 48962 34244 48974
rect 34300 49028 34356 49038
rect 34300 48934 34356 48972
rect 33068 48862 33070 48914
rect 33122 48862 33124 48914
rect 33068 48850 33124 48862
rect 32956 48804 33012 48814
rect 32956 48710 33012 48748
rect 33292 48804 33348 48814
rect 33348 48748 33460 48804
rect 33292 48710 33348 48748
rect 33068 48580 33124 48590
rect 33068 47570 33124 48524
rect 33068 47518 33070 47570
rect 33122 47518 33124 47570
rect 33068 47460 33124 47518
rect 33068 47394 33124 47404
rect 33404 47348 33460 48748
rect 33852 48802 33908 48814
rect 34412 48804 34468 49646
rect 33852 48750 33854 48802
rect 33906 48750 33908 48802
rect 33628 48244 33684 48254
rect 33852 48244 33908 48750
rect 33628 48242 33908 48244
rect 33628 48190 33630 48242
rect 33682 48190 33908 48242
rect 33628 48188 33908 48190
rect 34300 48802 34468 48804
rect 34300 48750 34414 48802
rect 34466 48750 34468 48802
rect 34300 48748 34468 48750
rect 33180 47346 33460 47348
rect 33180 47294 33406 47346
rect 33458 47294 33460 47346
rect 33180 47292 33460 47294
rect 33068 46676 33124 46686
rect 32844 46674 33124 46676
rect 32844 46622 33070 46674
rect 33122 46622 33124 46674
rect 32844 46620 33124 46622
rect 32844 46002 32900 46620
rect 33068 46610 33124 46620
rect 32844 45950 32846 46002
rect 32898 45950 32900 46002
rect 32844 45938 32900 45950
rect 32956 46116 33012 46126
rect 32732 45838 32734 45890
rect 32786 45838 32788 45890
rect 32732 45668 32788 45838
rect 32956 45890 33012 46060
rect 32956 45838 32958 45890
rect 33010 45838 33012 45890
rect 32956 45826 33012 45838
rect 33180 45780 33236 47292
rect 33404 47282 33460 47292
rect 33516 48020 33572 48030
rect 33516 46786 33572 47964
rect 33628 47012 33684 48188
rect 33852 47684 33908 47694
rect 33740 47460 33796 47470
rect 33740 47366 33796 47404
rect 33628 46946 33684 46956
rect 33740 47124 33796 47134
rect 33852 47124 33908 47628
rect 34188 47236 34244 47246
rect 34300 47236 34356 48748
rect 34412 48738 34468 48748
rect 34636 48804 34692 48814
rect 34636 48710 34692 48748
rect 34860 47684 34916 47694
rect 34860 47458 34916 47628
rect 34860 47406 34862 47458
rect 34914 47406 34916 47458
rect 34860 47394 34916 47406
rect 34636 47348 34692 47358
rect 34244 47180 34356 47236
rect 34412 47346 34692 47348
rect 34412 47294 34638 47346
rect 34690 47294 34692 47346
rect 34412 47292 34692 47294
rect 34188 47170 34244 47180
rect 33796 47068 33908 47124
rect 33516 46734 33518 46786
rect 33570 46734 33572 46786
rect 33516 46722 33572 46734
rect 33180 45686 33236 45724
rect 33292 46674 33348 46686
rect 33292 46622 33294 46674
rect 33346 46622 33348 46674
rect 33292 46452 33348 46622
rect 33740 46674 33796 47068
rect 34076 46900 34132 46910
rect 33740 46622 33742 46674
rect 33794 46622 33796 46674
rect 33740 46610 33796 46622
rect 33964 46844 34076 46900
rect 33964 46452 34020 46844
rect 34076 46806 34132 46844
rect 32732 45602 32788 45612
rect 33292 45556 33348 46396
rect 33628 46396 34020 46452
rect 33628 46114 33684 46396
rect 33628 46062 33630 46114
rect 33682 46062 33684 46114
rect 33628 46050 33684 46062
rect 33964 46004 34020 46014
rect 33964 46002 34244 46004
rect 33964 45950 33966 46002
rect 34018 45950 34244 46002
rect 33964 45948 34244 45950
rect 33964 45938 34020 45948
rect 32508 45014 32564 45052
rect 33180 45500 33348 45556
rect 33852 45666 33908 45678
rect 33852 45614 33854 45666
rect 33906 45614 33908 45666
rect 32396 44548 32452 44558
rect 32396 44324 32452 44492
rect 32396 44322 33012 44324
rect 32396 44270 32398 44322
rect 32450 44270 33012 44322
rect 32396 44268 33012 44270
rect 32396 44258 32452 44268
rect 32060 44100 32116 44110
rect 32060 43650 32116 44044
rect 32060 43598 32062 43650
rect 32114 43598 32116 43650
rect 32060 41972 32116 43598
rect 32508 43428 32564 43438
rect 32508 43334 32564 43372
rect 32060 41906 32116 41916
rect 32956 42642 33012 44268
rect 33180 43708 33236 45500
rect 33404 45108 33460 45118
rect 33404 45014 33460 45052
rect 33852 44548 33908 45614
rect 33852 44482 33908 44492
rect 33516 44436 33572 44446
rect 33516 44342 33572 44380
rect 33068 43652 33236 43708
rect 33292 44322 33348 44334
rect 33292 44270 33294 44322
rect 33346 44270 33348 44322
rect 33068 42868 33124 43652
rect 33068 42802 33124 42812
rect 33180 43538 33236 43550
rect 33180 43486 33182 43538
rect 33234 43486 33236 43538
rect 33180 43428 33236 43486
rect 33292 43540 33348 44270
rect 34188 44322 34244 45948
rect 34412 46002 34468 47292
rect 34636 47282 34692 47292
rect 34412 45950 34414 46002
rect 34466 45950 34468 46002
rect 34412 45938 34468 45950
rect 34524 46564 34580 46574
rect 34524 45890 34580 46508
rect 34524 45838 34526 45890
rect 34578 45838 34580 45890
rect 34524 45826 34580 45838
rect 34748 45780 34804 45790
rect 34748 45686 34804 45724
rect 34300 45668 34356 45678
rect 34300 45574 34356 45612
rect 34972 45332 35028 50318
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35532 49308 35700 49364
rect 35532 49138 35588 49308
rect 35644 49252 35700 49308
rect 35868 49252 35924 49262
rect 35644 49250 35924 49252
rect 35644 49198 35870 49250
rect 35922 49198 35924 49250
rect 35644 49196 35924 49198
rect 35868 49186 35924 49196
rect 35532 49086 35534 49138
rect 35586 49086 35588 49138
rect 35532 49074 35588 49086
rect 35084 49028 35140 49038
rect 35084 48934 35140 48972
rect 35420 49028 35476 49066
rect 35420 48962 35476 48972
rect 35980 49028 36036 52108
rect 35644 48914 35700 48926
rect 35644 48862 35646 48914
rect 35698 48862 35700 48914
rect 35644 48804 35700 48862
rect 35308 48748 35700 48804
rect 35980 48804 36036 48972
rect 36092 48804 36148 48814
rect 35980 48802 36148 48804
rect 35980 48750 36094 48802
rect 36146 48750 36148 48802
rect 35980 48748 36148 48750
rect 35308 48020 35364 48748
rect 35084 47964 35364 48020
rect 35644 48468 35700 48478
rect 35084 47460 35140 47964
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35644 47684 35700 48412
rect 35644 47570 35700 47628
rect 35644 47518 35646 47570
rect 35698 47518 35700 47570
rect 35196 47460 35252 47470
rect 35084 47458 35252 47460
rect 35084 47406 35198 47458
rect 35250 47406 35252 47458
rect 35084 47404 35252 47406
rect 35084 47234 35140 47246
rect 35084 47182 35086 47234
rect 35138 47182 35140 47234
rect 35084 46788 35140 47182
rect 35196 47124 35252 47404
rect 35196 47058 35252 47068
rect 35084 46722 35140 46732
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35644 45668 35700 47518
rect 35700 45612 35812 45668
rect 35644 45602 35700 45612
rect 35644 45332 35700 45342
rect 34188 44270 34190 44322
rect 34242 44270 34244 44322
rect 34188 44258 34244 44270
rect 34524 45276 35028 45332
rect 35532 45276 35644 45332
rect 34524 44546 34580 45276
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34524 44494 34526 44546
rect 34578 44494 34580 44546
rect 33964 43764 34020 43774
rect 33404 43652 33460 43662
rect 33404 43558 33460 43596
rect 33292 43474 33348 43484
rect 33964 43538 34020 43708
rect 33964 43486 33966 43538
rect 34018 43486 34020 43538
rect 33964 43474 34020 43486
rect 32956 42590 32958 42642
rect 33010 42590 33012 42642
rect 32172 41858 32228 41870
rect 32172 41806 32174 41858
rect 32226 41806 32228 41858
rect 32172 40852 32228 41806
rect 32956 41186 33012 42590
rect 33180 42194 33236 43372
rect 33516 43316 33572 43326
rect 33516 42754 33572 43260
rect 33852 42980 33908 42990
rect 33852 42866 33908 42924
rect 33852 42814 33854 42866
rect 33906 42814 33908 42866
rect 33852 42802 33908 42814
rect 33516 42702 33518 42754
rect 33570 42702 33572 42754
rect 33516 42690 33572 42702
rect 34524 42308 34580 44494
rect 35420 44436 35476 44446
rect 35532 44436 35588 45276
rect 35644 45266 35700 45276
rect 35420 44434 35588 44436
rect 35420 44382 35422 44434
rect 35474 44382 35588 44434
rect 35420 44380 35588 44382
rect 34748 44324 34804 44334
rect 34748 44230 34804 44268
rect 35420 44324 35476 44380
rect 35420 44258 35476 44268
rect 34972 44210 35028 44222
rect 34972 44158 34974 44210
rect 35026 44158 35028 44210
rect 34636 44098 34692 44110
rect 34636 44046 34638 44098
rect 34690 44046 34692 44098
rect 34636 43650 34692 44046
rect 34636 43598 34638 43650
rect 34690 43598 34692 43650
rect 34636 43586 34692 43598
rect 34972 43652 35028 44158
rect 34748 42868 34804 42878
rect 34748 42774 34804 42812
rect 34524 42242 34580 42252
rect 33180 42142 33182 42194
rect 33234 42142 33236 42194
rect 33180 42130 33236 42142
rect 34524 42082 34580 42094
rect 34524 42030 34526 42082
rect 34578 42030 34580 42082
rect 33964 41972 34020 41982
rect 32956 41134 32958 41186
rect 33010 41134 33012 41186
rect 32956 41122 33012 41134
rect 33852 41748 33908 41758
rect 33852 41186 33908 41692
rect 33852 41134 33854 41186
rect 33906 41134 33908 41186
rect 33852 41122 33908 41134
rect 32956 40964 33012 40974
rect 32956 40870 33012 40908
rect 32172 40786 32228 40796
rect 33964 40628 34020 41916
rect 34524 41972 34580 42030
rect 34300 41748 34356 41758
rect 34188 41746 34356 41748
rect 34188 41694 34302 41746
rect 34354 41694 34356 41746
rect 34188 41692 34356 41694
rect 34076 40628 34132 40638
rect 33964 40626 34132 40628
rect 33964 40574 34078 40626
rect 34130 40574 34132 40626
rect 33964 40572 34132 40574
rect 34076 40562 34132 40572
rect 32284 40404 32340 40414
rect 32284 39730 32340 40348
rect 32284 39678 32286 39730
rect 32338 39678 32340 39730
rect 32284 39666 32340 39678
rect 34076 39620 34132 39630
rect 34188 39620 34244 41692
rect 34300 41682 34356 41692
rect 34524 40852 34580 41916
rect 34972 42084 35028 43596
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35308 42868 35364 42878
rect 35084 42084 35140 42094
rect 34972 42082 35140 42084
rect 34972 42030 35086 42082
rect 35138 42030 35140 42082
rect 34972 42028 35140 42030
rect 34636 41748 34692 41758
rect 34636 41746 34804 41748
rect 34636 41694 34638 41746
rect 34690 41694 34804 41746
rect 34636 41692 34804 41694
rect 34636 41682 34692 41692
rect 34524 40626 34580 40796
rect 34524 40574 34526 40626
rect 34578 40574 34580 40626
rect 34524 40562 34580 40574
rect 34636 41188 34692 41198
rect 34636 40290 34692 41132
rect 34748 40404 34804 41692
rect 34860 41188 34916 41198
rect 34972 41188 35028 42028
rect 35084 42018 35140 42028
rect 35308 41970 35364 42812
rect 35308 41918 35310 41970
rect 35362 41918 35364 41970
rect 35308 41906 35364 41918
rect 35420 42308 35476 42318
rect 35420 41748 35476 42252
rect 35532 42194 35588 42206
rect 35532 42142 35534 42194
rect 35586 42142 35588 42194
rect 35532 41972 35588 42142
rect 35756 42196 35812 45612
rect 35980 42756 36036 48748
rect 36092 48738 36148 48748
rect 36316 48468 36372 52444
rect 36428 51268 36484 51278
rect 36876 51268 36932 54350
rect 37100 52948 37156 52958
rect 36988 52276 37044 52286
rect 36988 52182 37044 52220
rect 37100 52274 37156 52892
rect 37100 52222 37102 52274
rect 37154 52222 37156 52274
rect 37100 52210 37156 52222
rect 37212 52722 37268 52734
rect 37212 52670 37214 52722
rect 37266 52670 37268 52722
rect 37212 52164 37268 52670
rect 37324 52500 37380 55134
rect 37772 55074 37828 55086
rect 37772 55022 37774 55074
rect 37826 55022 37828 55074
rect 37660 53956 37716 53966
rect 37660 53844 37716 53900
rect 37772 53844 37828 55022
rect 38108 55074 38164 55086
rect 38108 55022 38110 55074
rect 38162 55022 38164 55074
rect 38108 54740 38164 55022
rect 38108 53956 38164 54684
rect 38220 54516 38276 54526
rect 38220 54422 38276 54460
rect 38108 53890 38164 53900
rect 38220 53844 38276 53854
rect 38332 53844 38388 55246
rect 40236 55298 40292 55310
rect 40236 55246 40238 55298
rect 40290 55246 40292 55298
rect 39004 55074 39060 55086
rect 39004 55022 39006 55074
rect 39058 55022 39060 55074
rect 38892 54626 38948 54638
rect 38892 54574 38894 54626
rect 38946 54574 38948 54626
rect 38556 54516 38612 54526
rect 38556 54422 38612 54460
rect 38892 54516 38948 54574
rect 38892 54450 38948 54460
rect 39004 54404 39060 55022
rect 39900 55076 39956 55086
rect 39900 54982 39956 55020
rect 40236 55076 40292 55246
rect 40236 55010 40292 55020
rect 41020 55186 41076 55198
rect 41020 55134 41022 55186
rect 41074 55134 41076 55186
rect 41020 54738 41076 55134
rect 41020 54686 41022 54738
rect 41074 54686 41076 54738
rect 41020 54674 41076 54686
rect 41916 55076 41972 55086
rect 39564 54628 39620 54638
rect 40908 54628 40964 54638
rect 39564 54534 39620 54572
rect 40796 54572 40908 54628
rect 39004 54338 39060 54348
rect 39228 54514 39284 54526
rect 39228 54462 39230 54514
rect 39282 54462 39284 54514
rect 37660 53842 38052 53844
rect 37660 53790 37662 53842
rect 37714 53790 38052 53842
rect 37660 53788 38052 53790
rect 37660 53778 37716 53788
rect 37996 53732 38052 53788
rect 38276 53788 38388 53844
rect 38780 54068 38836 54078
rect 38220 53732 38276 53788
rect 37996 53730 38276 53732
rect 37996 53678 38222 53730
rect 38274 53678 38276 53730
rect 37996 53676 38276 53678
rect 38220 53666 38276 53676
rect 37996 53508 38052 53518
rect 37996 53506 38164 53508
rect 37996 53454 37998 53506
rect 38050 53454 38164 53506
rect 37996 53452 38164 53454
rect 37996 53442 38052 53452
rect 37324 52434 37380 52444
rect 37212 52098 37268 52108
rect 37324 52162 37380 52174
rect 37324 52110 37326 52162
rect 37378 52110 37380 52162
rect 37324 51716 37380 52110
rect 37324 51650 37380 51660
rect 38108 51716 38164 53452
rect 38668 52388 38724 52398
rect 38668 52274 38724 52332
rect 38668 52222 38670 52274
rect 38722 52222 38724 52274
rect 38668 52210 38724 52222
rect 38220 52164 38276 52174
rect 38220 52070 38276 52108
rect 38108 51650 38164 51660
rect 36428 51266 36932 51268
rect 36428 51214 36430 51266
rect 36482 51214 36932 51266
rect 36428 51212 36932 51214
rect 37996 51604 38052 51614
rect 36428 50596 36484 51212
rect 37996 50706 38052 51548
rect 38780 51380 38836 54012
rect 38892 53844 38948 53854
rect 39228 53844 39284 54462
rect 40348 54404 40404 54414
rect 40348 54310 40404 54348
rect 38948 53788 39284 53844
rect 38892 53750 38948 53788
rect 40796 53060 40852 54572
rect 40908 54534 40964 54572
rect 41132 54514 41188 54526
rect 41132 54462 41134 54514
rect 41186 54462 41188 54514
rect 41132 54404 41188 54462
rect 41356 54516 41412 54526
rect 41356 54422 41412 54460
rect 41468 54514 41524 54526
rect 41468 54462 41470 54514
rect 41522 54462 41524 54514
rect 40908 53956 40964 53966
rect 40908 53862 40964 53900
rect 41132 53172 41188 54348
rect 41244 53956 41300 53966
rect 41468 53956 41524 54462
rect 41244 53954 41524 53956
rect 41244 53902 41246 53954
rect 41298 53902 41524 53954
rect 41244 53900 41524 53902
rect 41580 54516 41636 54526
rect 41244 53890 41300 53900
rect 41244 53732 41300 53742
rect 41244 53638 41300 53676
rect 41356 53172 41412 53182
rect 41132 53116 41300 53172
rect 40908 53060 40964 53070
rect 40796 53058 40964 53060
rect 40796 53006 40910 53058
rect 40962 53006 40964 53058
rect 40796 53004 40964 53006
rect 40348 52836 40404 52846
rect 40348 52742 40404 52780
rect 40236 52162 40292 52174
rect 40236 52110 40238 52162
rect 40290 52110 40292 52162
rect 39116 52052 39172 52062
rect 39116 51958 39172 51996
rect 38892 51604 38948 51642
rect 38892 51538 38948 51548
rect 40124 51604 40180 51614
rect 40124 51510 40180 51548
rect 39676 51492 39732 51502
rect 39676 51398 39732 51436
rect 40236 51492 40292 52110
rect 40348 51492 40404 51502
rect 40236 51490 40404 51492
rect 40236 51438 40350 51490
rect 40402 51438 40404 51490
rect 40236 51436 40404 51438
rect 39116 51380 39172 51390
rect 39452 51380 39508 51390
rect 38780 51324 38948 51380
rect 38556 51268 38612 51278
rect 38556 51174 38612 51212
rect 37996 50654 37998 50706
rect 38050 50654 38052 50706
rect 37996 50642 38052 50654
rect 36428 50502 36484 50540
rect 37324 50596 37380 50606
rect 37324 49810 37380 50540
rect 37324 49758 37326 49810
rect 37378 49758 37380 49810
rect 36540 49698 36596 49710
rect 36540 49646 36542 49698
rect 36594 49646 36596 49698
rect 36540 49250 36596 49646
rect 37324 49700 37380 49758
rect 38444 49924 38500 49934
rect 37772 49700 37828 49710
rect 37324 49698 37828 49700
rect 37324 49646 37774 49698
rect 37826 49646 37828 49698
rect 37324 49644 37828 49646
rect 37772 49588 37828 49644
rect 37772 49532 38276 49588
rect 36540 49198 36542 49250
rect 36594 49198 36596 49250
rect 36540 49186 36596 49198
rect 36316 48402 36372 48412
rect 38220 48132 38276 49532
rect 38444 49140 38500 49868
rect 38444 49138 38612 49140
rect 38444 49086 38446 49138
rect 38498 49086 38612 49138
rect 38444 49084 38612 49086
rect 38444 49074 38500 49084
rect 38556 48468 38612 49084
rect 38780 48468 38836 48478
rect 38220 48038 38276 48076
rect 38444 48466 38836 48468
rect 38444 48414 38782 48466
rect 38834 48414 38836 48466
rect 38444 48412 38836 48414
rect 38108 47460 38164 47470
rect 38108 47366 38164 47404
rect 38444 46898 38500 48412
rect 38780 48402 38836 48412
rect 38892 48356 38948 51324
rect 39116 51378 39396 51380
rect 39116 51326 39118 51378
rect 39170 51326 39396 51378
rect 39116 51324 39396 51326
rect 39116 51314 39172 51324
rect 39228 51156 39284 51166
rect 39340 51156 39396 51324
rect 39452 51286 39508 51324
rect 40012 51156 40068 51166
rect 39340 51154 40068 51156
rect 39340 51102 40014 51154
rect 40066 51102 40068 51154
rect 39340 51100 40068 51102
rect 39228 51062 39284 51100
rect 40012 51090 40068 51100
rect 40124 50708 40180 50718
rect 40236 50708 40292 51436
rect 40348 51426 40404 51436
rect 40908 51492 40964 53004
rect 41132 52946 41188 52958
rect 41132 52894 41134 52946
rect 41186 52894 41188 52946
rect 41132 52836 41188 52894
rect 41132 52770 41188 52780
rect 41244 52724 41300 53116
rect 41356 53078 41412 53116
rect 41468 52724 41524 52734
rect 41580 52724 41636 54460
rect 41692 53844 41748 53854
rect 41692 52946 41748 53788
rect 41692 52894 41694 52946
rect 41746 52894 41748 52946
rect 41692 52882 41748 52894
rect 41916 52948 41972 55020
rect 42028 53844 42084 53854
rect 42028 53750 42084 53788
rect 42924 53732 42980 55356
rect 43148 55346 43204 55356
rect 43596 55076 43652 55086
rect 43708 55076 43764 56030
rect 45500 55412 45556 59200
rect 47740 56308 47796 59200
rect 47740 56242 47796 56252
rect 48972 56308 49028 56318
rect 48972 56214 49028 56252
rect 49980 56308 50036 59200
rect 52220 57428 52276 59200
rect 52220 57372 52388 57428
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49980 56242 50036 56252
rect 52220 56308 52276 56318
rect 52220 56214 52276 56252
rect 47740 56084 47796 56094
rect 47964 56084 48020 56094
rect 47740 56082 48020 56084
rect 47740 56030 47742 56082
rect 47794 56030 47966 56082
rect 48018 56030 48020 56082
rect 47740 56028 48020 56030
rect 45500 55346 45556 55356
rect 46732 55412 46788 55422
rect 46732 55318 46788 55356
rect 45724 55298 45780 55310
rect 45724 55246 45726 55298
rect 45778 55246 45780 55298
rect 43484 55074 43764 55076
rect 43484 55022 43598 55074
rect 43650 55022 43764 55074
rect 43484 55020 43764 55022
rect 45388 55076 45444 55086
rect 45724 55076 45780 55246
rect 45388 55074 45780 55076
rect 45388 55022 45390 55074
rect 45442 55022 45780 55074
rect 45388 55020 45780 55022
rect 43484 54068 43540 55020
rect 43596 54982 43652 55020
rect 43484 54002 43540 54012
rect 42364 53620 42420 53630
rect 42364 53618 42644 53620
rect 42364 53566 42366 53618
rect 42418 53566 42644 53618
rect 42364 53564 42644 53566
rect 42364 53554 42420 53564
rect 42140 53508 42196 53518
rect 42140 53506 42308 53508
rect 42140 53454 42142 53506
rect 42194 53454 42308 53506
rect 42140 53452 42308 53454
rect 42140 53442 42196 53452
rect 42028 52948 42084 52958
rect 41916 52946 42084 52948
rect 41916 52894 42030 52946
rect 42082 52894 42084 52946
rect 41916 52892 42084 52894
rect 41244 52668 41412 52724
rect 41244 52500 41300 52510
rect 41244 52274 41300 52444
rect 41244 52222 41246 52274
rect 41298 52222 41300 52274
rect 41020 51492 41076 51502
rect 40964 51490 41076 51492
rect 40964 51438 41022 51490
rect 41074 51438 41076 51490
rect 40964 51436 41076 51438
rect 40908 51398 40964 51436
rect 41020 51426 41076 51436
rect 41244 51490 41300 52222
rect 41244 51438 41246 51490
rect 41298 51438 41300 51490
rect 41244 51426 41300 51438
rect 40124 50706 40292 50708
rect 40124 50654 40126 50706
rect 40178 50654 40292 50706
rect 40124 50652 40292 50654
rect 40348 51268 40404 51278
rect 40124 50642 40180 50652
rect 38892 48290 38948 48300
rect 39116 48356 39172 48366
rect 39116 48354 39284 48356
rect 39116 48302 39118 48354
rect 39170 48302 39284 48354
rect 39116 48300 39284 48302
rect 39116 48290 39172 48300
rect 38556 47460 38612 47470
rect 38556 47366 38612 47404
rect 39004 47458 39060 47470
rect 39004 47406 39006 47458
rect 39058 47406 39060 47458
rect 38780 47236 38836 47246
rect 39004 47236 39060 47406
rect 38780 47234 39060 47236
rect 38780 47182 38782 47234
rect 38834 47182 39060 47234
rect 38780 47180 39060 47182
rect 38780 47170 38836 47180
rect 38444 46846 38446 46898
rect 38498 46846 38500 46898
rect 36652 46788 36708 46798
rect 36652 46694 36708 46732
rect 37324 46674 37380 46686
rect 37324 46622 37326 46674
rect 37378 46622 37380 46674
rect 37100 44996 37156 45006
rect 37324 44996 37380 46622
rect 38444 46564 38500 46846
rect 38780 47012 38836 47022
rect 38780 46786 38836 46956
rect 38780 46734 38782 46786
rect 38834 46734 38836 46786
rect 38780 46722 38836 46734
rect 38444 46498 38500 46508
rect 38668 46450 38724 46462
rect 38668 46398 38670 46450
rect 38722 46398 38724 46450
rect 38668 45892 38724 46398
rect 38668 45826 38724 45836
rect 38668 45668 38724 45678
rect 38668 45574 38724 45612
rect 37100 44994 37380 44996
rect 37100 44942 37102 44994
rect 37154 44942 37380 44994
rect 37100 44940 37380 44942
rect 36204 44548 36260 44558
rect 36204 43708 36260 44492
rect 37100 44324 37156 44940
rect 37100 43764 37156 44268
rect 36204 43652 36484 43708
rect 35980 42690 36036 42700
rect 35756 42140 36260 42196
rect 35532 41906 35588 41916
rect 35868 41972 35924 41982
rect 35868 41970 36148 41972
rect 35868 41918 35870 41970
rect 35922 41918 36148 41970
rect 35868 41916 36148 41918
rect 35868 41906 35924 41916
rect 35532 41748 35588 41758
rect 35420 41746 35700 41748
rect 35420 41694 35534 41746
rect 35586 41694 35700 41746
rect 35420 41692 35700 41694
rect 35532 41682 35588 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35420 41412 35476 41422
rect 35644 41412 35700 41692
rect 35308 41410 35700 41412
rect 35308 41358 35422 41410
rect 35474 41358 35700 41410
rect 35308 41356 35700 41358
rect 34860 41186 35028 41188
rect 34860 41134 34862 41186
rect 34914 41134 35028 41186
rect 34860 41132 35028 41134
rect 34860 41122 34916 41132
rect 34972 40514 35028 41132
rect 35196 41186 35252 41198
rect 35196 41134 35198 41186
rect 35250 41134 35252 41186
rect 35196 41076 35252 41134
rect 35196 41010 35252 41020
rect 35308 40964 35364 41356
rect 35420 41346 35476 41356
rect 36092 41298 36148 41916
rect 36204 41412 36260 42140
rect 36316 41860 36372 41870
rect 36316 41766 36372 41804
rect 36204 41356 36372 41412
rect 36092 41246 36094 41298
rect 36146 41246 36148 41298
rect 36092 41234 36148 41246
rect 35420 41188 35476 41198
rect 35420 41094 35476 41132
rect 35980 41074 36036 41086
rect 35980 41022 35982 41074
rect 36034 41022 36036 41074
rect 35644 40964 35700 40974
rect 35308 40908 35476 40964
rect 34972 40462 34974 40514
rect 35026 40462 35028 40514
rect 34972 40450 35028 40462
rect 35308 40628 35364 40638
rect 34748 40338 34804 40348
rect 35308 40402 35364 40572
rect 35308 40350 35310 40402
rect 35362 40350 35364 40402
rect 35308 40338 35364 40350
rect 35420 40402 35476 40908
rect 35644 40962 35924 40964
rect 35644 40910 35646 40962
rect 35698 40910 35924 40962
rect 35644 40908 35924 40910
rect 35644 40898 35700 40908
rect 35756 40626 35812 40638
rect 35756 40574 35758 40626
rect 35810 40574 35812 40626
rect 35420 40350 35422 40402
rect 35474 40350 35476 40402
rect 35420 40338 35476 40350
rect 35532 40404 35588 40414
rect 35532 40310 35588 40348
rect 34636 40238 34638 40290
rect 34690 40238 34692 40290
rect 34636 40226 34692 40238
rect 34300 40178 34356 40190
rect 34300 40126 34302 40178
rect 34354 40126 34356 40178
rect 34300 39732 34356 40126
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34300 39676 34916 39732
rect 34076 39618 34244 39620
rect 34076 39566 34078 39618
rect 34130 39566 34244 39618
rect 34076 39564 34244 39566
rect 34860 39620 34916 39676
rect 34972 39620 35028 39630
rect 34860 39618 35028 39620
rect 34860 39566 34974 39618
rect 35026 39566 35028 39618
rect 34860 39564 35028 39566
rect 34076 39554 34132 39564
rect 33852 39508 33908 39518
rect 33516 39506 33908 39508
rect 33516 39454 33854 39506
rect 33906 39454 33908 39506
rect 33516 39452 33908 39454
rect 31948 38770 32004 38780
rect 32396 38946 32452 38958
rect 32396 38894 32398 38946
rect 32450 38894 32452 38946
rect 32396 38668 32452 38894
rect 31836 37998 31838 38050
rect 31890 37998 31892 38050
rect 31836 37986 31892 37998
rect 32284 38612 32452 38668
rect 32508 38834 32564 38846
rect 32508 38782 32510 38834
rect 32562 38782 32564 38834
rect 32508 38612 32564 38782
rect 32060 37940 32116 37950
rect 32060 37846 32116 37884
rect 32172 37938 32228 37950
rect 32172 37886 32174 37938
rect 32226 37886 32228 37938
rect 31724 37762 31780 37772
rect 32172 37828 32228 37886
rect 32172 37762 32228 37772
rect 32284 37604 32340 38612
rect 32508 38546 32564 38556
rect 32956 38612 33012 38622
rect 31276 37214 31278 37266
rect 31330 37214 31332 37266
rect 31276 37202 31332 37214
rect 31388 37548 31556 37604
rect 32060 37548 32340 37604
rect 32396 38500 32452 38510
rect 31388 35364 31444 37548
rect 32060 37492 32116 37548
rect 31500 37490 32116 37492
rect 31500 37438 32062 37490
rect 32114 37438 32116 37490
rect 31500 37436 32116 37438
rect 31500 37380 31556 37436
rect 31500 37266 31556 37324
rect 31500 37214 31502 37266
rect 31554 37214 31556 37266
rect 31500 37202 31556 37214
rect 31724 36594 31780 37436
rect 32060 37426 32116 37436
rect 32284 37380 32340 37390
rect 32396 37380 32452 38444
rect 32956 38162 33012 38556
rect 33516 38612 33572 39452
rect 33852 39442 33908 39452
rect 33628 38836 33684 38846
rect 33628 38668 33684 38780
rect 33852 38724 33908 38734
rect 33628 38612 33796 38668
rect 33852 38630 33908 38668
rect 33516 38546 33572 38556
rect 32956 38110 32958 38162
rect 33010 38110 33012 38162
rect 32956 38098 33012 38110
rect 33404 38050 33460 38062
rect 33404 37998 33406 38050
rect 33458 37998 33460 38050
rect 33404 37940 33460 37998
rect 33292 37828 33348 37838
rect 32956 37492 33012 37502
rect 32284 37378 32452 37380
rect 32284 37326 32286 37378
rect 32338 37326 32452 37378
rect 32284 37324 32452 37326
rect 32284 37314 32340 37324
rect 32060 37268 32116 37278
rect 31948 37156 32004 37166
rect 31948 37062 32004 37100
rect 31724 36542 31726 36594
rect 31778 36542 31780 36594
rect 31724 36530 31780 36542
rect 31388 35298 31444 35308
rect 31724 35700 31780 35710
rect 31724 34804 31780 35644
rect 31724 34738 31780 34748
rect 31836 34690 31892 34702
rect 31836 34638 31838 34690
rect 31890 34638 31892 34690
rect 31388 34130 31444 34142
rect 31388 34078 31390 34130
rect 31442 34078 31444 34130
rect 31388 33124 31444 34078
rect 31388 33058 31444 33068
rect 31500 30210 31556 30222
rect 31500 30158 31502 30210
rect 31554 30158 31556 30210
rect 31500 30100 31556 30158
rect 31500 30034 31556 30044
rect 31836 29204 31892 34638
rect 32060 31892 32116 37212
rect 32396 37268 32452 37324
rect 32396 37202 32452 37212
rect 32844 37436 32956 37492
rect 32172 36482 32228 36494
rect 32172 36430 32174 36482
rect 32226 36430 32228 36482
rect 32172 34916 32228 36430
rect 32844 36482 32900 37436
rect 32956 37426 33012 37436
rect 32844 36430 32846 36482
rect 32898 36430 32900 36482
rect 32844 35700 32900 36430
rect 33292 36594 33348 37772
rect 33292 36542 33294 36594
rect 33346 36542 33348 36594
rect 33068 35700 33124 35710
rect 32620 35698 33124 35700
rect 32620 35646 33070 35698
rect 33122 35646 33124 35698
rect 32620 35644 33124 35646
rect 32396 34916 32452 34926
rect 32172 34850 32228 34860
rect 32284 34914 32452 34916
rect 32284 34862 32398 34914
rect 32450 34862 32452 34914
rect 32284 34860 32452 34862
rect 32284 33460 32340 34860
rect 32396 34850 32452 34860
rect 32508 34130 32564 34142
rect 32508 34078 32510 34130
rect 32562 34078 32564 34130
rect 32396 33906 32452 33918
rect 32396 33854 32398 33906
rect 32450 33854 32452 33906
rect 32396 33796 32452 33854
rect 32508 33908 32564 34078
rect 32508 33842 32564 33852
rect 32396 33730 32452 33740
rect 32396 33460 32452 33470
rect 32284 33404 32396 33460
rect 32396 33394 32452 33404
rect 32620 33346 32676 35644
rect 33068 35634 33124 35644
rect 33292 35476 33348 36542
rect 32956 35420 33348 35476
rect 32732 34916 32788 34926
rect 32956 34916 33012 35420
rect 33180 35252 33236 35262
rect 32732 34914 33012 34916
rect 32732 34862 32734 34914
rect 32786 34862 33012 34914
rect 32732 34860 33012 34862
rect 33068 34916 33124 34926
rect 32732 34850 32788 34860
rect 32620 33294 32622 33346
rect 32674 33294 32676 33346
rect 32620 33282 32676 33294
rect 33068 33796 33124 34860
rect 33180 34802 33236 35196
rect 33180 34750 33182 34802
rect 33234 34750 33236 34802
rect 33180 34738 33236 34750
rect 33068 32562 33124 33740
rect 33404 33460 33460 37884
rect 33516 36036 33572 36046
rect 33516 35364 33572 35980
rect 33516 35298 33572 35308
rect 33628 34020 33684 34030
rect 33740 34020 33796 38612
rect 34188 38164 34244 39564
rect 34748 39506 34804 39518
rect 34748 39454 34750 39506
rect 34802 39454 34804 39506
rect 34300 38948 34356 38958
rect 34748 38948 34804 39454
rect 34300 38946 34804 38948
rect 34300 38894 34302 38946
rect 34354 38894 34804 38946
rect 34300 38892 34804 38894
rect 34300 38668 34356 38892
rect 34972 38834 35028 39564
rect 35644 39060 35700 39070
rect 35532 39004 35644 39060
rect 35532 38946 35588 39004
rect 35644 38994 35700 39004
rect 35532 38894 35534 38946
rect 35586 38894 35588 38946
rect 35532 38882 35588 38894
rect 35756 38948 35812 40574
rect 35756 38882 35812 38892
rect 34972 38782 34974 38834
rect 35026 38782 35028 38834
rect 34300 38612 34468 38668
rect 34300 38164 34356 38174
rect 34244 38162 34356 38164
rect 34244 38110 34302 38162
rect 34354 38110 34356 38162
rect 34244 38108 34356 38110
rect 34188 38070 34244 38108
rect 34300 38098 34356 38108
rect 33852 37828 33908 37838
rect 33852 37734 33908 37772
rect 34412 37492 34468 38612
rect 33964 37436 34468 37492
rect 33964 34468 34020 37436
rect 34300 37268 34356 37278
rect 34076 36258 34132 36270
rect 34076 36206 34078 36258
rect 34130 36206 34132 36258
rect 34076 35700 34132 36206
rect 34076 35634 34132 35644
rect 34188 35586 34244 35598
rect 34188 35534 34190 35586
rect 34242 35534 34244 35586
rect 34188 35364 34244 35534
rect 34188 35298 34244 35308
rect 34300 34804 34356 37212
rect 34860 37266 34916 37278
rect 34860 37214 34862 37266
rect 34914 37214 34916 37266
rect 34636 36596 34692 36606
rect 34636 36502 34692 36540
rect 34748 35924 34804 35934
rect 34748 35830 34804 35868
rect 34860 35812 34916 37214
rect 34860 35746 34916 35756
rect 34748 35698 34804 35710
rect 34748 35646 34750 35698
rect 34802 35646 34804 35698
rect 34748 35364 34804 35646
rect 34524 34804 34580 34814
rect 34300 34802 34580 34804
rect 34300 34750 34526 34802
rect 34578 34750 34580 34802
rect 34300 34748 34580 34750
rect 34524 34738 34580 34748
rect 34636 34692 34692 34702
rect 34636 34598 34692 34636
rect 33964 34412 34132 34468
rect 33628 34018 33796 34020
rect 33628 33966 33630 34018
rect 33682 33966 33796 34018
rect 33628 33964 33796 33966
rect 33964 34242 34020 34254
rect 33964 34190 33966 34242
rect 34018 34190 34020 34242
rect 33628 33954 33684 33964
rect 33404 33394 33460 33404
rect 33516 33572 33572 33582
rect 33516 33458 33572 33516
rect 33516 33406 33518 33458
rect 33570 33406 33572 33458
rect 33516 33394 33572 33406
rect 33628 32676 33684 32686
rect 33068 32510 33070 32562
rect 33122 32510 33124 32562
rect 32060 31826 32116 31836
rect 32396 31892 32452 31902
rect 32396 31554 32452 31836
rect 33068 31892 33124 32510
rect 33068 31826 33124 31836
rect 33404 32620 33628 32676
rect 33404 31666 33460 32620
rect 33628 32582 33684 32620
rect 33964 32676 34020 34190
rect 33964 32610 34020 32620
rect 33404 31614 33406 31666
rect 33458 31614 33460 31666
rect 33404 31602 33460 31614
rect 33964 31778 34020 31790
rect 33964 31726 33966 31778
rect 34018 31726 34020 31778
rect 32396 31502 32398 31554
rect 32450 31502 32452 31554
rect 32396 31490 32452 31502
rect 33180 31220 33236 31230
rect 33180 31126 33236 31164
rect 33964 30996 34020 31726
rect 33964 30930 34020 30940
rect 34076 31108 34132 34412
rect 34748 34356 34804 35308
rect 34972 34468 35028 38782
rect 35532 38724 35588 38734
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35308 37268 35364 37278
rect 35532 37268 35588 38668
rect 35868 37380 35924 40908
rect 35980 38668 36036 41022
rect 36204 40962 36260 40974
rect 36204 40910 36206 40962
rect 36258 40910 36260 40962
rect 36204 40852 36260 40910
rect 36204 40786 36260 40796
rect 36316 40628 36372 41356
rect 36316 40534 36372 40572
rect 36428 39060 36484 43652
rect 36988 43652 37156 43708
rect 37212 44434 37268 44446
rect 37212 44382 37214 44434
rect 37266 44382 37268 44434
rect 37212 43652 37268 44382
rect 36764 43426 36820 43438
rect 36764 43374 36766 43426
rect 36818 43374 36820 43426
rect 36764 40516 36820 43374
rect 36764 40450 36820 40460
rect 36876 42756 36932 42766
rect 36876 41076 36932 42700
rect 36764 40292 36820 40302
rect 36876 40292 36932 41020
rect 36764 40290 36932 40292
rect 36764 40238 36766 40290
rect 36818 40238 36932 40290
rect 36764 40236 36932 40238
rect 36988 41186 37044 43652
rect 37212 43586 37268 43596
rect 37436 44212 37492 44222
rect 37436 43650 37492 44156
rect 37436 43598 37438 43650
rect 37490 43598 37492 43650
rect 37436 43586 37492 43598
rect 38780 43652 38836 43662
rect 38892 43652 38948 47180
rect 39116 46674 39172 46686
rect 39116 46622 39118 46674
rect 39170 46622 39172 46674
rect 39116 46564 39172 46622
rect 39116 46498 39172 46508
rect 39228 46676 39284 48300
rect 39676 48132 39732 48142
rect 39676 48038 39732 48076
rect 40012 47572 40068 47582
rect 39452 47570 40068 47572
rect 39452 47518 40014 47570
rect 40066 47518 40068 47570
rect 39452 47516 40068 47518
rect 39452 47234 39508 47516
rect 40012 47506 40068 47516
rect 39452 47182 39454 47234
rect 39506 47182 39508 47234
rect 39452 47012 39508 47182
rect 39452 46946 39508 46956
rect 39564 47234 39620 47246
rect 39564 47182 39566 47234
rect 39618 47182 39620 47234
rect 39228 45892 39284 46620
rect 39452 46786 39508 46798
rect 39452 46734 39454 46786
rect 39506 46734 39508 46786
rect 39452 46564 39508 46734
rect 39564 46788 39620 47182
rect 39564 46722 39620 46732
rect 39676 47234 39732 47246
rect 39676 47182 39678 47234
rect 39730 47182 39732 47234
rect 39676 46564 39732 47182
rect 40348 47012 40404 51212
rect 41132 51266 41188 51278
rect 41132 51214 41134 51266
rect 41186 51214 41188 51266
rect 40908 50596 40964 50606
rect 40908 50502 40964 50540
rect 41132 50484 41188 51214
rect 41356 50820 41412 52668
rect 41468 52722 41636 52724
rect 41468 52670 41470 52722
rect 41522 52670 41636 52722
rect 41468 52668 41636 52670
rect 41468 51378 41524 52668
rect 41468 51326 41470 51378
rect 41522 51326 41524 51378
rect 41468 51156 41524 51326
rect 41468 51090 41524 51100
rect 41692 51940 41748 51950
rect 41916 51940 41972 52892
rect 42028 52882 42084 52892
rect 42140 52052 42196 52062
rect 42140 51958 42196 51996
rect 41692 51938 41972 51940
rect 41692 51886 41694 51938
rect 41746 51886 41972 51938
rect 41692 51884 41972 51886
rect 41132 50418 41188 50428
rect 41244 50764 41412 50820
rect 40348 46956 41188 47012
rect 40348 46898 40404 46956
rect 40348 46846 40350 46898
rect 40402 46846 40404 46898
rect 40348 46834 40404 46846
rect 40908 46788 40964 46798
rect 40908 46694 40964 46732
rect 41132 46786 41188 46956
rect 41132 46734 41134 46786
rect 41186 46734 41188 46786
rect 41132 46722 41188 46734
rect 39452 46508 39732 46564
rect 39004 45836 39284 45892
rect 39004 45218 39060 45836
rect 39228 45668 39284 45678
rect 39284 45612 39396 45668
rect 39228 45602 39284 45612
rect 39004 45166 39006 45218
rect 39058 45166 39060 45218
rect 39004 45154 39060 45166
rect 39228 45330 39284 45342
rect 39228 45278 39230 45330
rect 39282 45278 39284 45330
rect 39228 44436 39284 45278
rect 39340 45218 39396 45612
rect 39340 45166 39342 45218
rect 39394 45166 39396 45218
rect 39340 45154 39396 45166
rect 39564 45106 39620 45118
rect 39564 45054 39566 45106
rect 39618 45054 39620 45106
rect 39340 44436 39396 44446
rect 39228 44434 39396 44436
rect 39228 44382 39342 44434
rect 39394 44382 39396 44434
rect 39228 44380 39396 44382
rect 39340 44370 39396 44380
rect 39564 43762 39620 45054
rect 39564 43710 39566 43762
rect 39618 43710 39620 43762
rect 39564 43698 39620 43710
rect 39676 43764 39732 46508
rect 40236 46676 40292 46686
rect 40012 44324 40068 44334
rect 40012 44230 40068 44268
rect 39228 43652 39284 43662
rect 38892 43650 39284 43652
rect 38892 43598 39230 43650
rect 39282 43598 39284 43650
rect 38892 43596 39284 43598
rect 38780 43558 38836 43596
rect 37324 43540 37380 43550
rect 37324 43446 37380 43484
rect 39228 43540 39284 43596
rect 39452 43652 39508 43662
rect 39452 43558 39508 43596
rect 39676 43650 39732 43708
rect 39676 43598 39678 43650
rect 39730 43598 39732 43650
rect 39676 43586 39732 43598
rect 39228 43474 39284 43484
rect 38668 43316 38724 43326
rect 38668 43222 38724 43260
rect 40124 42756 40180 42766
rect 40236 42756 40292 46620
rect 41244 46564 41300 50764
rect 41356 50596 41412 50606
rect 41692 50596 41748 51884
rect 42252 51604 42308 53452
rect 42588 52836 42644 53564
rect 42812 53172 42868 53182
rect 42812 53058 42868 53116
rect 42812 53006 42814 53058
rect 42866 53006 42868 53058
rect 42812 52994 42868 53006
rect 42588 52274 42644 52780
rect 42588 52222 42590 52274
rect 42642 52222 42644 52274
rect 42588 52210 42644 52222
rect 42252 51510 42308 51548
rect 42476 52162 42532 52174
rect 42476 52110 42478 52162
rect 42530 52110 42532 52162
rect 41804 51378 41860 51390
rect 41804 51326 41806 51378
rect 41858 51326 41860 51378
rect 41804 51268 41860 51326
rect 42140 51268 42196 51278
rect 41804 51266 42196 51268
rect 41804 51214 42142 51266
rect 42194 51214 42196 51266
rect 41804 51212 42196 51214
rect 42140 51202 42196 51212
rect 42476 51154 42532 52110
rect 42924 52162 42980 53676
rect 42924 52110 42926 52162
rect 42978 52110 42980 52162
rect 42924 52098 42980 52110
rect 44604 53844 44660 53854
rect 42476 51102 42478 51154
rect 42530 51102 42532 51154
rect 42476 50708 42532 51102
rect 42476 50642 42532 50652
rect 44156 50708 44212 50718
rect 44156 50614 44212 50652
rect 41412 50540 41748 50596
rect 41356 50502 41412 50540
rect 42028 50484 42084 50494
rect 42028 50390 42084 50428
rect 42812 48132 42868 48142
rect 42812 47458 42868 48076
rect 42812 47406 42814 47458
rect 42866 47406 42868 47458
rect 42812 47394 42868 47406
rect 41356 47348 41412 47358
rect 41356 46898 41412 47292
rect 42140 47348 42196 47358
rect 42140 47254 42196 47292
rect 41356 46846 41358 46898
rect 41410 46846 41412 46898
rect 41356 46834 41412 46846
rect 41468 46676 41524 46686
rect 41524 46620 41972 46676
rect 41468 46582 41524 46620
rect 41020 46508 41300 46564
rect 41020 46002 41076 46508
rect 41020 45950 41022 46002
rect 41074 45950 41076 46002
rect 41020 45332 41076 45950
rect 41244 46004 41300 46508
rect 41244 45948 41636 46004
rect 41580 45890 41636 45948
rect 41580 45838 41582 45890
rect 41634 45838 41636 45890
rect 41580 45826 41636 45838
rect 41916 45890 41972 46620
rect 41916 45838 41918 45890
rect 41970 45838 41972 45890
rect 41916 45826 41972 45838
rect 41356 45780 41412 45790
rect 41020 45266 41076 45276
rect 41132 45778 41412 45780
rect 41132 45726 41358 45778
rect 41410 45726 41412 45778
rect 41132 45724 41412 45726
rect 41020 44996 41076 45006
rect 40572 44322 40628 44334
rect 40572 44270 40574 44322
rect 40626 44270 40628 44322
rect 40572 43652 40628 44270
rect 40572 43586 40628 43596
rect 40908 44324 40964 44334
rect 40348 42756 40404 42766
rect 40236 42754 40404 42756
rect 40236 42702 40350 42754
rect 40402 42702 40404 42754
rect 40236 42700 40404 42702
rect 40124 42662 40180 42700
rect 40348 42690 40404 42700
rect 40684 42756 40740 42794
rect 40684 42690 40740 42700
rect 40684 42530 40740 42542
rect 40684 42478 40686 42530
rect 40738 42478 40740 42530
rect 37772 41972 37828 41982
rect 37772 41298 37828 41916
rect 40124 41860 40180 41870
rect 40124 41766 40180 41804
rect 40012 41748 40068 41758
rect 40684 41748 40740 42478
rect 40908 41970 40964 44268
rect 41020 44322 41076 44940
rect 41132 44434 41188 45724
rect 41356 45714 41412 45724
rect 41804 45666 41860 45678
rect 41804 45614 41806 45666
rect 41858 45614 41860 45666
rect 41804 45332 41860 45614
rect 41804 45276 42420 45332
rect 42364 45218 42420 45276
rect 42364 45166 42366 45218
rect 42418 45166 42420 45218
rect 42364 45154 42420 45166
rect 41132 44382 41134 44434
rect 41186 44382 41188 44434
rect 41132 44370 41188 44382
rect 41580 45106 41636 45118
rect 41580 45054 41582 45106
rect 41634 45054 41636 45106
rect 41020 44270 41022 44322
rect 41074 44270 41076 44322
rect 41020 44212 41076 44270
rect 41580 44324 41636 45054
rect 44492 44996 44548 45006
rect 44492 44902 44548 44940
rect 41580 44258 41636 44268
rect 41020 44146 41076 44156
rect 41244 44098 41300 44110
rect 41244 44046 41246 44098
rect 41298 44046 41300 44098
rect 41132 43764 41188 43802
rect 41244 43764 41300 44046
rect 41188 43708 41300 43764
rect 41132 43698 41188 43708
rect 41580 43652 41636 43662
rect 41580 43558 41636 43596
rect 41356 43538 41412 43550
rect 41356 43486 41358 43538
rect 41410 43486 41412 43538
rect 41244 43428 41300 43438
rect 41020 43426 41300 43428
rect 41020 43374 41246 43426
rect 41298 43374 41300 43426
rect 41020 43372 41300 43374
rect 41020 42754 41076 43372
rect 41244 43362 41300 43372
rect 41020 42702 41022 42754
rect 41074 42702 41076 42754
rect 41020 42690 41076 42702
rect 40908 41918 40910 41970
rect 40962 41918 40964 41970
rect 40908 41906 40964 41918
rect 41356 41972 41412 43486
rect 44604 42980 44660 53788
rect 44940 52836 44996 52846
rect 44940 52742 44996 52780
rect 45388 49028 45444 55020
rect 45388 48962 45444 48972
rect 47740 47572 47796 56028
rect 47964 56018 48020 56028
rect 51212 56082 51268 56094
rect 51212 56030 51214 56082
rect 51266 56030 51268 56082
rect 51212 55468 51268 56030
rect 50876 55412 51268 55468
rect 52332 55412 52388 57372
rect 54460 56308 54516 59200
rect 54460 56242 54516 56252
rect 56028 56308 56084 56318
rect 56028 56214 56084 56252
rect 54572 56084 54628 56094
rect 55020 56084 55076 56094
rect 54572 56082 55076 56084
rect 54572 56030 54574 56082
rect 54626 56030 55022 56082
rect 55074 56030 55076 56082
rect 54572 56028 55076 56030
rect 50876 55074 50932 55412
rect 52332 55346 52388 55356
rect 53676 55412 53732 55422
rect 53676 55318 53732 55356
rect 52668 55298 52724 55310
rect 52668 55246 52670 55298
rect 52722 55246 52724 55298
rect 50876 55022 50878 55074
rect 50930 55022 50932 55074
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50876 53844 50932 55022
rect 52108 55076 52164 55086
rect 52668 55076 52724 55246
rect 52108 55074 52724 55076
rect 52108 55022 52110 55074
rect 52162 55022 52724 55074
rect 52108 55020 52724 55022
rect 52108 55010 52164 55020
rect 47740 47506 47796 47516
rect 50316 53788 50932 53844
rect 50316 46004 50372 53788
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50316 45938 50372 45948
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 44604 42914 44660 42924
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 41356 41906 41412 41916
rect 41692 41858 41748 41870
rect 41692 41806 41694 41858
rect 41746 41806 41748 41858
rect 41692 41748 41748 41806
rect 43820 41860 43876 41870
rect 43820 41766 43876 41804
rect 40684 41692 41748 41748
rect 40012 41654 40068 41692
rect 37772 41246 37774 41298
rect 37826 41246 37828 41298
rect 37772 41234 37828 41246
rect 39900 41298 39956 41310
rect 39900 41246 39902 41298
rect 39954 41246 39956 41298
rect 36988 41134 36990 41186
rect 37042 41134 37044 41186
rect 36764 40226 36820 40236
rect 36428 38668 36484 39004
rect 36876 38836 36932 38846
rect 36764 38834 36932 38836
rect 36764 38782 36878 38834
rect 36930 38782 36932 38834
rect 36764 38780 36932 38782
rect 35980 38612 36148 38668
rect 36428 38612 36708 38668
rect 35980 37380 36036 37390
rect 35868 37378 36036 37380
rect 35868 37326 35982 37378
rect 36034 37326 36036 37378
rect 35868 37324 36036 37326
rect 35980 37314 36036 37324
rect 35308 37266 35588 37268
rect 35308 37214 35310 37266
rect 35362 37214 35588 37266
rect 35308 37212 35588 37214
rect 36092 37268 36148 38612
rect 35308 37202 35364 37212
rect 36092 37202 36148 37212
rect 36316 36932 36372 36942
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 36092 36596 36148 36606
rect 35420 36370 35476 36382
rect 35420 36318 35422 36370
rect 35474 36318 35476 36370
rect 35420 36036 35476 36318
rect 35532 36036 35588 36046
rect 35420 35980 35532 36036
rect 35588 35980 35700 36036
rect 35532 35970 35588 35980
rect 35644 35810 35700 35980
rect 35644 35758 35646 35810
rect 35698 35758 35700 35810
rect 35644 35746 35700 35758
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 34916 35140 34926
rect 35084 34822 35140 34860
rect 36092 34802 36148 36540
rect 36316 36484 36372 36876
rect 36652 36708 36708 38612
rect 36764 36932 36820 38780
rect 36876 38770 36932 38780
rect 36988 38724 37044 41134
rect 38444 40516 38500 40526
rect 38220 38948 38276 38958
rect 38220 38854 38276 38892
rect 36988 38658 37044 38668
rect 37436 38834 37492 38846
rect 37436 38782 37438 38834
rect 37490 38782 37492 38834
rect 37436 38724 37492 38782
rect 37436 38658 37492 38668
rect 37772 38724 37828 38734
rect 37212 38276 37268 38286
rect 37212 38162 37268 38220
rect 37212 38110 37214 38162
rect 37266 38110 37268 38162
rect 37212 38098 37268 38110
rect 37772 38052 37828 38668
rect 37772 38050 37940 38052
rect 37772 37998 37774 38050
rect 37826 37998 37940 38050
rect 37772 37996 37940 37998
rect 37772 37986 37828 37996
rect 36764 36866 36820 36876
rect 36652 36652 37044 36708
rect 36652 36596 36708 36652
rect 36652 36530 36708 36540
rect 36988 36594 37044 36652
rect 36988 36542 36990 36594
rect 37042 36542 37044 36594
rect 36988 36530 37044 36542
rect 36204 34916 36260 34926
rect 36316 34916 36372 36428
rect 37548 36258 37604 36270
rect 37548 36206 37550 36258
rect 37602 36206 37604 36258
rect 37324 35812 37380 35822
rect 37380 35756 37492 35812
rect 37324 35746 37380 35756
rect 36428 35586 36484 35598
rect 36428 35534 36430 35586
rect 36482 35534 36484 35586
rect 36428 35364 36484 35534
rect 36428 35298 36484 35308
rect 36204 34914 36372 34916
rect 36204 34862 36206 34914
rect 36258 34862 36372 34914
rect 36204 34860 36372 34862
rect 37324 34914 37380 34926
rect 37324 34862 37326 34914
rect 37378 34862 37380 34914
rect 36204 34850 36260 34860
rect 36092 34750 36094 34802
rect 36146 34750 36148 34802
rect 36092 34738 36148 34750
rect 34972 34402 35028 34412
rect 36316 34580 36372 34590
rect 34636 34300 34804 34356
rect 34412 34132 34468 34142
rect 34412 34038 34468 34076
rect 34300 33572 34356 33582
rect 34188 33460 34244 33470
rect 34188 31108 34244 33404
rect 34300 31778 34356 33516
rect 34636 33348 34692 34300
rect 34860 34244 34916 34254
rect 34860 34242 35364 34244
rect 34860 34190 34862 34242
rect 34914 34190 35364 34242
rect 34860 34188 35364 34190
rect 34860 34178 34916 34188
rect 34748 34130 34804 34142
rect 34748 34078 34750 34130
rect 34802 34078 34804 34130
rect 34748 33572 34804 34078
rect 35308 34132 35364 34188
rect 35308 34076 35588 34132
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34804 33516 35140 33572
rect 34748 33506 34804 33516
rect 34748 33348 34804 33358
rect 34300 31726 34302 31778
rect 34354 31726 34356 31778
rect 34300 31714 34356 31726
rect 34524 33346 34804 33348
rect 34524 33294 34750 33346
rect 34802 33294 34804 33346
rect 34524 33292 34804 33294
rect 34524 31780 34580 33292
rect 34748 33282 34804 33292
rect 34860 33234 34916 33246
rect 34860 33182 34862 33234
rect 34914 33182 34916 33234
rect 34860 32676 34916 33182
rect 34524 31714 34580 31724
rect 34636 32620 34916 32676
rect 34300 31108 34356 31118
rect 34188 31106 34356 31108
rect 34188 31054 34302 31106
rect 34354 31054 34356 31106
rect 34188 31052 34356 31054
rect 31948 30212 32004 30222
rect 31948 30118 32004 30156
rect 34076 29540 34132 31052
rect 34300 30324 34356 31052
rect 34412 30324 34468 30334
rect 34300 30322 34468 30324
rect 34300 30270 34414 30322
rect 34466 30270 34468 30322
rect 34300 30268 34468 30270
rect 34412 30258 34468 30268
rect 34636 30212 34692 32620
rect 35084 32564 35140 33516
rect 35308 33124 35364 33134
rect 35308 33030 35364 33068
rect 35532 32676 35588 34076
rect 35868 33908 35924 33918
rect 35868 33346 35924 33852
rect 35868 33294 35870 33346
rect 35922 33294 35924 33346
rect 35868 33282 35924 33294
rect 36316 33234 36372 34524
rect 37324 34356 37380 34862
rect 37436 34802 37492 35756
rect 37548 35364 37604 36206
rect 37660 36036 37716 36046
rect 37660 35922 37716 35980
rect 37660 35870 37662 35922
rect 37714 35870 37716 35922
rect 37660 35858 37716 35870
rect 37772 35812 37828 35822
rect 37772 35718 37828 35756
rect 37548 35298 37604 35308
rect 37436 34750 37438 34802
rect 37490 34750 37492 34802
rect 37436 34580 37492 34750
rect 37548 34804 37604 34814
rect 37548 34690 37604 34748
rect 37548 34638 37550 34690
rect 37602 34638 37604 34690
rect 37548 34626 37604 34638
rect 37436 34514 37492 34524
rect 36988 34300 37828 34356
rect 36652 34132 36708 34142
rect 36652 34038 36708 34076
rect 36316 33182 36318 33234
rect 36370 33182 36372 33234
rect 36316 33170 36372 33182
rect 36204 32676 36260 32686
rect 35532 32674 36260 32676
rect 35532 32622 36206 32674
rect 36258 32622 36260 32674
rect 35532 32620 36260 32622
rect 34972 32562 35140 32564
rect 34972 32510 35086 32562
rect 35138 32510 35140 32562
rect 34972 32508 35140 32510
rect 34860 32452 34916 32462
rect 34636 30146 34692 30156
rect 34748 32450 34916 32452
rect 34748 32398 34862 32450
rect 34914 32398 34916 32450
rect 34748 32396 34916 32398
rect 34748 29764 34804 32396
rect 34860 32386 34916 32396
rect 34860 30996 34916 31006
rect 34972 30996 35028 32508
rect 35084 32498 35140 32508
rect 35756 32452 35812 32462
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35756 31108 35812 32396
rect 36092 31668 36148 31678
rect 36204 31668 36260 32620
rect 36988 32004 37044 34300
rect 37772 34242 37828 34300
rect 37772 34190 37774 34242
rect 37826 34190 37828 34242
rect 37772 34178 37828 34190
rect 37100 34130 37156 34142
rect 37100 34078 37102 34130
rect 37154 34078 37156 34130
rect 37100 33908 37156 34078
rect 37100 33842 37156 33852
rect 37100 33348 37156 33358
rect 37100 33254 37156 33292
rect 37772 33348 37828 33358
rect 37884 33348 37940 37996
rect 37996 38050 38052 38062
rect 37996 37998 37998 38050
rect 38050 37998 38052 38050
rect 37996 37156 38052 37998
rect 38220 38050 38276 38062
rect 38220 37998 38222 38050
rect 38274 37998 38276 38050
rect 38220 37492 38276 37998
rect 38220 37426 38276 37436
rect 38444 37938 38500 40460
rect 39900 38724 39956 41246
rect 52668 40964 52724 55020
rect 54572 53844 54628 56028
rect 55020 56018 55076 56028
rect 56700 55410 56756 59200
rect 56700 55358 56702 55410
rect 56754 55358 56756 55410
rect 56700 55346 56756 55358
rect 55580 55298 55636 55310
rect 55580 55246 55582 55298
rect 55634 55246 55636 55298
rect 55244 54404 55300 54414
rect 55580 54404 55636 55246
rect 55244 54402 55636 54404
rect 55244 54350 55246 54402
rect 55298 54350 55636 54402
rect 55244 54348 55636 54350
rect 55244 54338 55300 54348
rect 54572 53778 54628 53788
rect 55356 44436 55412 54348
rect 55356 44370 55412 44380
rect 52668 40898 52724 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 39900 38658 39956 38668
rect 40348 38722 40404 38734
rect 40348 38670 40350 38722
rect 40402 38670 40404 38722
rect 38444 37886 38446 37938
rect 38498 37886 38500 37938
rect 38108 37156 38164 37166
rect 37996 37154 38164 37156
rect 37996 37102 38110 37154
rect 38162 37102 38164 37154
rect 37996 37100 38164 37102
rect 38108 35924 38164 37100
rect 38108 35698 38164 35868
rect 38108 35646 38110 35698
rect 38162 35646 38164 35698
rect 38108 35634 38164 35646
rect 37828 33292 37940 33348
rect 38220 34356 38276 34366
rect 38444 34356 38500 37886
rect 39564 37492 39620 37502
rect 39564 37398 39620 37436
rect 39900 37492 39956 37502
rect 40348 37492 40404 38670
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 39900 37490 40404 37492
rect 39900 37438 39902 37490
rect 39954 37438 40404 37490
rect 39900 37436 40404 37438
rect 39900 37426 39956 37436
rect 40348 37378 40404 37436
rect 40348 37326 40350 37378
rect 40402 37326 40404 37378
rect 40348 37314 40404 37326
rect 40236 37042 40292 37054
rect 40236 36990 40238 37042
rect 40290 36990 40292 37042
rect 38892 36594 38948 36606
rect 38892 36542 38894 36594
rect 38946 36542 38948 36594
rect 38892 36484 38948 36542
rect 38276 34300 38500 34356
rect 38668 35924 38724 35934
rect 37772 33282 37828 33292
rect 37212 33124 37268 33134
rect 37212 33030 37268 33068
rect 37548 32452 37604 32462
rect 37548 32358 37604 32396
rect 36148 31612 36260 31668
rect 36876 31948 37044 32004
rect 36092 31574 36148 31612
rect 35756 31014 35812 31052
rect 34860 30994 35028 30996
rect 34860 30942 34862 30994
rect 34914 30942 35028 30994
rect 34860 30940 35028 30942
rect 35980 30996 36036 31006
rect 34860 30930 34916 30940
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34860 30212 34916 30222
rect 34860 30118 34916 30156
rect 35868 30212 35924 30222
rect 35868 30118 35924 30156
rect 34748 29708 34916 29764
rect 34188 29540 34244 29550
rect 34076 29538 34244 29540
rect 34076 29486 34190 29538
rect 34242 29486 34244 29538
rect 34076 29484 34244 29486
rect 34188 29474 34244 29484
rect 31836 29138 31892 29148
rect 31164 28130 31220 28140
rect 29932 28084 29988 28094
rect 29932 27990 29988 28028
rect 30828 28084 30884 28094
rect 30828 27990 30884 28028
rect 30268 27972 30324 27982
rect 30268 27878 30324 27916
rect 29372 27806 29374 27858
rect 29426 27806 29428 27858
rect 29260 27524 29316 27534
rect 28252 26404 28308 26414
rect 28252 25618 28308 26348
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28252 25554 28308 25566
rect 29260 25618 29316 27468
rect 29260 25566 29262 25618
rect 29314 25566 29316 25618
rect 29260 25508 29316 25566
rect 29260 25442 29316 25452
rect 29372 25172 29428 27806
rect 34860 25620 34916 29708
rect 35644 29650 35700 29662
rect 35644 29598 35646 29650
rect 35698 29598 35700 29650
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35644 28084 35700 29598
rect 35868 29428 35924 29438
rect 35980 29428 36036 30940
rect 36876 30996 36932 31948
rect 36988 31780 37044 31790
rect 36988 31686 37044 31724
rect 37884 31780 37940 31790
rect 36876 30902 36932 30940
rect 37100 31666 37156 31678
rect 37100 31614 37102 31666
rect 37154 31614 37156 31666
rect 36204 30324 36260 30334
rect 36204 30230 36260 30268
rect 36988 30212 37044 30222
rect 37100 30212 37156 31614
rect 37324 31668 37380 31678
rect 37212 31556 37268 31566
rect 37212 31462 37268 31500
rect 37044 30156 37156 30212
rect 37324 30882 37380 31612
rect 37324 30830 37326 30882
rect 37378 30830 37380 30882
rect 36988 30146 37044 30156
rect 37324 29538 37380 30830
rect 37324 29486 37326 29538
rect 37378 29486 37380 29538
rect 37324 29474 37380 29486
rect 35868 29426 36036 29428
rect 35868 29374 35870 29426
rect 35922 29374 36036 29426
rect 35868 29372 36036 29374
rect 37884 29426 37940 31724
rect 38220 30994 38276 34300
rect 38668 34130 38724 35868
rect 38892 34916 38948 36428
rect 39564 36484 39620 36494
rect 40236 36484 40292 36990
rect 39564 36482 40292 36484
rect 39564 36430 39566 36482
rect 39618 36430 40292 36482
rect 39564 36428 40292 36430
rect 39340 35924 39396 35934
rect 39340 35830 39396 35868
rect 39340 34916 39396 34926
rect 38892 34914 39396 34916
rect 38892 34862 39342 34914
rect 39394 34862 39396 34914
rect 38892 34860 39396 34862
rect 39340 34850 39396 34860
rect 39228 34356 39284 34366
rect 39228 34262 39284 34300
rect 38668 34078 38670 34130
rect 38722 34078 38724 34130
rect 38668 34066 38724 34078
rect 39340 34244 39396 34254
rect 39340 33908 39396 34188
rect 39228 33852 39396 33908
rect 39228 33346 39284 33852
rect 39228 33294 39230 33346
rect 39282 33294 39284 33346
rect 39228 33282 39284 33294
rect 39564 33346 39620 36428
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 39788 35586 39844 35598
rect 39788 35534 39790 35586
rect 39842 35534 39844 35586
rect 39788 34244 39844 35534
rect 39788 34178 39844 34188
rect 39900 35364 39956 35374
rect 39900 34802 39956 35308
rect 39900 34750 39902 34802
rect 39954 34750 39956 34802
rect 39788 34018 39844 34030
rect 39788 33966 39790 34018
rect 39842 33966 39844 34018
rect 39788 33908 39844 33966
rect 39900 33908 39956 34750
rect 41916 35026 41972 35038
rect 41916 34974 41918 35026
rect 41970 34974 41972 35026
rect 41468 34690 41524 34702
rect 41468 34638 41470 34690
rect 41522 34638 41524 34690
rect 39788 33852 40180 33908
rect 39564 33294 39566 33346
rect 39618 33294 39620 33346
rect 39564 33282 39620 33294
rect 40012 33572 40068 33582
rect 38668 33236 38724 33246
rect 38444 33234 38724 33236
rect 38444 33182 38670 33234
rect 38722 33182 38724 33234
rect 38444 33180 38724 33182
rect 38332 33124 38388 33134
rect 38444 33124 38500 33180
rect 38668 33170 38724 33180
rect 38388 33068 38500 33124
rect 38332 33058 38388 33068
rect 38444 32562 38500 33068
rect 38444 32510 38446 32562
rect 38498 32510 38500 32562
rect 38444 32498 38500 32510
rect 39004 33122 39060 33134
rect 39004 33070 39006 33122
rect 39058 33070 39060 33122
rect 38220 30942 38222 30994
rect 38274 30942 38276 30994
rect 38220 30324 38276 30942
rect 38220 30258 38276 30268
rect 37884 29374 37886 29426
rect 37938 29374 37940 29426
rect 35868 29362 35924 29372
rect 37884 29362 37940 29374
rect 35644 28018 35700 28028
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34860 25554 34916 25564
rect 29372 25106 29428 25116
rect 39004 24612 39060 33070
rect 39564 32676 39620 32686
rect 39564 32450 39620 32620
rect 40012 32562 40068 33516
rect 40124 33234 40180 33852
rect 41468 33572 41524 34638
rect 41916 34580 41972 34974
rect 41916 34514 41972 34524
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 41468 33506 41524 33516
rect 40124 33182 40126 33234
rect 40178 33182 40180 33234
rect 40124 33170 40180 33182
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 40012 32510 40014 32562
rect 40066 32510 40068 32562
rect 40012 32498 40068 32510
rect 39564 32398 39566 32450
rect 39618 32398 39620 32450
rect 39564 31948 39620 32398
rect 39564 31892 39732 31948
rect 39116 31780 39172 31790
rect 39116 31686 39172 31724
rect 39676 31666 39732 31892
rect 39676 31614 39678 31666
rect 39730 31614 39732 31666
rect 39676 31602 39732 31614
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 39004 24546 39060 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 19068 22866 19124 22876
rect 28028 22866 28084 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 6748 9650 6804 9660
rect 5628 9426 5684 9436
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 5068 6738 5124 6748
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 2492 4226 2548 4238
rect 2492 4174 2494 4226
rect 2546 4174 2548 4226
rect 2492 3892 2548 4174
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 2492 3826 2548 3836
rect 2268 3666 2436 3668
rect 2268 3614 2270 3666
rect 2322 3614 2436 3666
rect 2268 3612 2436 3614
rect 2268 3602 2324 3612
rect 1708 3442 1764 3454
rect 1708 3390 1710 3442
rect 1762 3390 1764 3442
rect 1708 3332 1764 3390
rect 1708 2100 1764 3276
rect 2716 3442 2772 3454
rect 2716 3390 2718 3442
rect 2770 3390 2772 3442
rect 2716 3332 2772 3390
rect 2716 3266 2772 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 1708 2034 1764 2044
<< via2 >>
rect 2156 57596 2212 57652
rect 1708 55804 1764 55860
rect 2156 56028 2212 56084
rect 1596 54572 1652 54628
rect 1484 44828 1540 44884
rect 924 42252 980 42308
rect 1036 39564 1092 39620
rect 1372 36204 1428 36260
rect 1036 32844 1092 32900
rect 1148 35644 1204 35700
rect 924 28700 980 28756
rect 1036 32396 1092 32452
rect 1148 23436 1204 23492
rect 1708 54012 1764 54068
rect 1708 52780 1764 52836
rect 1708 52220 1764 52276
rect 1820 51212 1876 51268
rect 1708 50706 1764 50708
rect 1708 50654 1710 50706
rect 1710 50654 1762 50706
rect 1762 50654 1764 50706
rect 1708 50652 1764 50654
rect 1708 50428 1764 50484
rect 2044 54626 2100 54628
rect 2044 54574 2046 54626
rect 2046 54574 2098 54626
rect 2098 54574 2100 54626
rect 2044 54572 2100 54574
rect 2044 51490 2100 51492
rect 2044 51438 2046 51490
rect 2046 51438 2098 51490
rect 2098 51438 2100 51490
rect 2044 51436 2100 51438
rect 2044 50652 2100 50708
rect 2268 49980 2324 50036
rect 1708 48636 1764 48692
rect 1708 46844 1764 46900
rect 1708 45276 1764 45332
rect 1708 45052 1764 45108
rect 2156 47628 2212 47684
rect 1820 43596 1876 43652
rect 1820 43260 1876 43316
rect 1708 41468 1764 41524
rect 1708 40236 1764 40292
rect 1708 39676 1764 39732
rect 2044 43484 2100 43540
rect 2268 44492 2324 44548
rect 2604 56082 2660 56084
rect 2604 56030 2606 56082
rect 2606 56030 2658 56082
rect 2658 56030 2660 56082
rect 2604 56028 2660 56030
rect 2492 54012 2548 54068
rect 3164 55804 3220 55860
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 5852 55132 5908 55188
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 2940 53788 2996 53844
rect 5628 53788 5684 53844
rect 2492 52834 2548 52836
rect 2492 52782 2494 52834
rect 2494 52782 2546 52834
rect 2546 52782 2548 52834
rect 2492 52780 2548 52782
rect 2492 51266 2548 51268
rect 2492 51214 2494 51266
rect 2494 51214 2546 51266
rect 2546 51214 2548 51266
rect 2492 51212 2548 51214
rect 2492 48636 2548 48692
rect 2492 46898 2548 46900
rect 2492 46846 2494 46898
rect 2494 46846 2546 46898
rect 2546 46846 2548 46898
rect 2492 46844 2548 46846
rect 2492 45276 2548 45332
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 3836 51884 3892 51940
rect 2716 51436 2772 51492
rect 2716 49980 2772 50036
rect 2716 48412 2772 48468
rect 2716 47458 2772 47460
rect 2716 47406 2718 47458
rect 2718 47406 2770 47458
rect 2770 47406 2772 47458
rect 2716 47404 2772 47406
rect 7980 53058 8036 53060
rect 7980 53006 7982 53058
rect 7982 53006 8034 53058
rect 8034 53006 8036 53058
rect 7980 53004 8036 53006
rect 5628 51436 5684 51492
rect 4396 51378 4452 51380
rect 4396 51326 4398 51378
rect 4398 51326 4450 51378
rect 4450 51326 4452 51378
rect 4396 51324 4452 51326
rect 5180 51324 5236 51380
rect 5068 51266 5124 51268
rect 5068 51214 5070 51266
rect 5070 51214 5122 51266
rect 5122 51214 5124 51266
rect 5068 51212 5124 51214
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 7644 51378 7700 51380
rect 7644 51326 7646 51378
rect 7646 51326 7698 51378
rect 7698 51326 7700 51378
rect 7644 51324 7700 51326
rect 5852 50764 5908 50820
rect 3836 49922 3892 49924
rect 3836 49870 3838 49922
rect 3838 49870 3890 49922
rect 3890 49870 3892 49922
rect 3836 49868 3892 49870
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 3052 48412 3108 48468
rect 3500 48466 3556 48468
rect 3500 48414 3502 48466
rect 3502 48414 3554 48466
rect 3554 48414 3556 48466
rect 3500 48412 3556 48414
rect 3276 47682 3332 47684
rect 3276 47630 3278 47682
rect 3278 47630 3330 47682
rect 3330 47630 3332 47682
rect 3276 47628 3332 47630
rect 3948 47458 4004 47460
rect 3948 47406 3950 47458
rect 3950 47406 4002 47458
rect 4002 47406 4004 47458
rect 3948 47404 4004 47406
rect 2268 42082 2324 42084
rect 2268 42030 2270 42082
rect 2270 42030 2322 42082
rect 2322 42030 2324 42082
rect 2268 42028 2324 42030
rect 2044 41916 2100 41972
rect 2716 43538 2772 43540
rect 2716 43486 2718 43538
rect 2718 43486 2770 43538
rect 2770 43486 2772 43538
rect 2716 43484 2772 43486
rect 2716 42642 2772 42644
rect 2716 42590 2718 42642
rect 2718 42590 2770 42642
rect 2770 42590 2772 42642
rect 2716 42588 2772 42590
rect 2044 39564 2100 39620
rect 1708 37938 1764 37940
rect 1708 37886 1710 37938
rect 1710 37886 1762 37938
rect 1762 37886 1764 37938
rect 1708 37884 1764 37886
rect 2044 37826 2100 37828
rect 2044 37774 2046 37826
rect 2046 37774 2098 37826
rect 2098 37774 2100 37826
rect 2044 37772 2100 37774
rect 1596 36428 1652 36484
rect 1708 37100 1764 37156
rect 1708 36092 1764 36148
rect 1484 28252 1540 28308
rect 1596 34412 1652 34468
rect 1372 15708 1428 15764
rect 1036 5852 1092 5908
rect 1708 34354 1764 34356
rect 1708 34302 1710 34354
rect 1710 34302 1762 34354
rect 1762 34302 1764 34354
rect 1708 34300 1764 34302
rect 1708 33234 1764 33236
rect 1708 33182 1710 33234
rect 1710 33182 1762 33234
rect 1762 33182 1764 33234
rect 1708 33180 1764 33182
rect 1708 32508 1764 32564
rect 2044 36540 2100 36596
rect 1932 36370 1988 36372
rect 1932 36318 1934 36370
rect 1934 36318 1986 36370
rect 1986 36318 1988 36370
rect 1932 36316 1988 36318
rect 1820 31052 1876 31108
rect 1932 35980 1988 36036
rect 1708 30716 1764 30772
rect 1708 27692 1764 27748
rect 1708 27132 1764 27188
rect 1708 25394 1764 25396
rect 1708 25342 1710 25394
rect 1710 25342 1762 25394
rect 1762 25342 1764 25394
rect 1708 25340 1764 25342
rect 2716 41970 2772 41972
rect 2716 41918 2718 41970
rect 2718 41918 2770 41970
rect 2770 41918 2772 41970
rect 2716 41916 2772 41918
rect 3164 44882 3220 44884
rect 3164 44830 3166 44882
rect 3166 44830 3218 44882
rect 3218 44830 3220 44882
rect 3164 44828 3220 44830
rect 3052 42530 3108 42532
rect 3052 42478 3054 42530
rect 3054 42478 3106 42530
rect 3106 42478 3108 42530
rect 3052 42476 3108 42478
rect 2492 40236 2548 40292
rect 2828 40236 2884 40292
rect 2940 39788 2996 39844
rect 3052 39618 3108 39620
rect 3052 39566 3054 39618
rect 3054 39566 3106 39618
rect 3106 39566 3108 39618
rect 3052 39564 3108 39566
rect 2604 39004 2660 39060
rect 2380 37660 2436 37716
rect 2044 35196 2100 35252
rect 2828 37826 2884 37828
rect 2828 37774 2830 37826
rect 2830 37774 2882 37826
rect 2882 37774 2884 37826
rect 2828 37772 2884 37774
rect 2604 37490 2660 37492
rect 2604 37438 2606 37490
rect 2606 37438 2658 37490
rect 2658 37438 2660 37490
rect 2604 37436 2660 37438
rect 2604 37042 2660 37044
rect 2604 36990 2606 37042
rect 2606 36990 2658 37042
rect 2658 36990 2660 37042
rect 2604 36988 2660 36990
rect 2940 36316 2996 36372
rect 2716 35980 2772 36036
rect 2940 35980 2996 36036
rect 2604 35922 2660 35924
rect 2604 35870 2606 35922
rect 2606 35870 2658 35922
rect 2658 35870 2660 35922
rect 2604 35868 2660 35870
rect 2716 35698 2772 35700
rect 2716 35646 2718 35698
rect 2718 35646 2770 35698
rect 2770 35646 2772 35698
rect 2716 35644 2772 35646
rect 2380 34972 2436 35028
rect 2940 35644 2996 35700
rect 2716 35196 2772 35252
rect 3164 37154 3220 37156
rect 3164 37102 3166 37154
rect 3166 37102 3218 37154
rect 3218 37102 3220 37154
rect 3164 37100 3220 37102
rect 3724 47068 3780 47124
rect 6076 48130 6132 48132
rect 6076 48078 6078 48130
rect 6078 48078 6130 48130
rect 6130 48078 6132 48130
rect 6076 48076 6132 48078
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4060 47068 4116 47124
rect 4508 46844 4564 46900
rect 4844 46786 4900 46788
rect 4844 46734 4846 46786
rect 4846 46734 4898 46786
rect 4898 46734 4900 46786
rect 4844 46732 4900 46734
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4508 45778 4564 45780
rect 4508 45726 4510 45778
rect 4510 45726 4562 45778
rect 4562 45726 4564 45778
rect 4508 45724 4564 45726
rect 4172 45388 4228 45444
rect 3724 44994 3780 44996
rect 3724 44942 3726 44994
rect 3726 44942 3778 44994
rect 3778 44942 3780 44994
rect 3724 44940 3780 44942
rect 3612 43596 3668 43652
rect 3388 40236 3444 40292
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4844 43596 4900 43652
rect 5292 43650 5348 43652
rect 5292 43598 5294 43650
rect 5294 43598 5346 43650
rect 5346 43598 5348 43650
rect 5292 43596 5348 43598
rect 4060 42140 4116 42196
rect 4060 41858 4116 41860
rect 4060 41806 4062 41858
rect 4062 41806 4114 41858
rect 4114 41806 4116 41858
rect 4060 41804 4116 41806
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5852 43426 5908 43428
rect 5852 43374 5854 43426
rect 5854 43374 5906 43426
rect 5906 43374 5908 43426
rect 5852 43372 5908 43374
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4284 40236 4340 40292
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5180 40460 5236 40516
rect 5068 40348 5124 40404
rect 4956 39900 5012 39956
rect 3388 39506 3444 39508
rect 3388 39454 3390 39506
rect 3390 39454 3442 39506
rect 3442 39454 3444 39506
rect 3388 39452 3444 39454
rect 3500 39394 3556 39396
rect 3500 39342 3502 39394
rect 3502 39342 3554 39394
rect 3554 39342 3556 39394
rect 3500 39340 3556 39342
rect 3836 39116 3892 39172
rect 3612 39004 3668 39060
rect 3500 38946 3556 38948
rect 3500 38894 3502 38946
rect 3502 38894 3554 38946
rect 3554 38894 3556 38946
rect 3500 38892 3556 38894
rect 3948 38780 4004 38836
rect 4172 39788 4228 39844
rect 4060 38556 4116 38612
rect 5740 40402 5796 40404
rect 5740 40350 5742 40402
rect 5742 40350 5794 40402
rect 5794 40350 5796 40402
rect 5740 40348 5796 40350
rect 5292 40236 5348 40292
rect 4284 39116 4340 39172
rect 4956 39116 5012 39172
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 5180 38834 5236 38836
rect 5180 38782 5182 38834
rect 5182 38782 5234 38834
rect 5234 38782 5236 38834
rect 5180 38780 5236 38782
rect 5628 39452 5684 39508
rect 5740 39058 5796 39060
rect 5740 39006 5742 39058
rect 5742 39006 5794 39058
rect 5794 39006 5796 39058
rect 5740 39004 5796 39006
rect 5628 38946 5684 38948
rect 5628 38894 5630 38946
rect 5630 38894 5682 38946
rect 5682 38894 5684 38946
rect 5628 38892 5684 38894
rect 6412 47852 6468 47908
rect 6636 48242 6692 48244
rect 6636 48190 6638 48242
rect 6638 48190 6690 48242
rect 6690 48190 6692 48242
rect 6636 48188 6692 48190
rect 7308 50818 7364 50820
rect 7308 50766 7310 50818
rect 7310 50766 7362 50818
rect 7362 50766 7364 50818
rect 7308 50764 7364 50766
rect 7084 48188 7140 48244
rect 6188 45500 6244 45556
rect 6524 45388 6580 45444
rect 6524 44716 6580 44772
rect 6188 43650 6244 43652
rect 6188 43598 6190 43650
rect 6190 43598 6242 43650
rect 6242 43598 6244 43650
rect 6188 43596 6244 43598
rect 7532 47404 7588 47460
rect 7308 47068 7364 47124
rect 7420 46620 7476 46676
rect 7420 46060 7476 46116
rect 6748 45388 6804 45444
rect 7084 45612 7140 45668
rect 6300 42252 6356 42308
rect 6412 42082 6468 42084
rect 6412 42030 6414 42082
rect 6414 42030 6466 42082
rect 6466 42030 6468 42082
rect 6412 42028 6468 42030
rect 6188 40514 6244 40516
rect 6188 40462 6190 40514
rect 6190 40462 6242 40514
rect 6242 40462 6244 40514
rect 6188 40460 6244 40462
rect 6188 40236 6244 40292
rect 6076 39900 6132 39956
rect 6860 44156 6916 44212
rect 6972 45500 7028 45556
rect 7196 44716 7252 44772
rect 6860 43372 6916 43428
rect 6636 43148 6692 43204
rect 6524 38834 6580 38836
rect 6524 38782 6526 38834
rect 6526 38782 6578 38834
rect 6578 38782 6580 38834
rect 6524 38780 6580 38782
rect 5292 38332 5348 38388
rect 4732 38050 4788 38052
rect 4732 37998 4734 38050
rect 4734 37998 4786 38050
rect 4786 37998 4788 38050
rect 4732 37996 4788 37998
rect 3612 37212 3668 37268
rect 3276 35980 3332 36036
rect 3836 36370 3892 36372
rect 3836 36318 3838 36370
rect 3838 36318 3890 36370
rect 3890 36318 3892 36370
rect 3836 36316 3892 36318
rect 3276 35698 3332 35700
rect 3276 35646 3278 35698
rect 3278 35646 3330 35698
rect 3330 35646 3332 35698
rect 3276 35644 3332 35646
rect 3052 35308 3108 35364
rect 2044 34748 2100 34804
rect 2940 34636 2996 34692
rect 2492 34524 2548 34580
rect 2492 34354 2548 34356
rect 2492 34302 2494 34354
rect 2494 34302 2546 34354
rect 2546 34302 2548 34354
rect 2492 34300 2548 34302
rect 2044 34242 2100 34244
rect 2044 34190 2046 34242
rect 2046 34190 2098 34242
rect 2098 34190 2100 34242
rect 2044 34188 2100 34190
rect 2044 33122 2100 33124
rect 2044 33070 2046 33122
rect 2046 33070 2098 33122
rect 2098 33070 2100 33122
rect 2044 33068 2100 33070
rect 2492 33234 2548 33236
rect 2492 33182 2494 33234
rect 2494 33182 2546 33234
rect 2546 33182 2548 33234
rect 2492 33180 2548 33182
rect 3164 34636 3220 34692
rect 3276 35252 3332 35308
rect 3052 33516 3108 33572
rect 2268 31836 2324 31892
rect 2156 30994 2212 30996
rect 2156 30942 2158 30994
rect 2158 30942 2210 30994
rect 2210 30942 2212 30994
rect 2156 30940 2212 30942
rect 2044 30268 2100 30324
rect 3836 35474 3892 35476
rect 3836 35422 3838 35474
rect 3838 35422 3890 35474
rect 3890 35422 3892 35474
rect 3836 35420 3892 35422
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4620 36428 4676 36484
rect 4060 35644 4116 35700
rect 3724 33404 3780 33460
rect 2828 32732 2884 32788
rect 3612 32562 3668 32564
rect 3612 32510 3614 32562
rect 3614 32510 3666 32562
rect 3666 32510 3668 32562
rect 3612 32508 3668 32510
rect 2380 29932 2436 29988
rect 2380 28924 2436 28980
rect 2268 28812 2324 28868
rect 2268 28642 2324 28644
rect 2268 28590 2270 28642
rect 2270 28590 2322 28642
rect 2322 28590 2324 28642
rect 2268 28588 2324 28590
rect 2044 28476 2100 28532
rect 2268 28364 2324 28420
rect 2156 27244 2212 27300
rect 2044 23826 2100 23828
rect 2044 23774 2046 23826
rect 2046 23774 2098 23826
rect 2098 23774 2100 23826
rect 2044 23772 2100 23774
rect 1708 23548 1764 23604
rect 1820 23436 1876 23492
rect 1708 21756 1764 21812
rect 3052 31778 3108 31780
rect 3052 31726 3054 31778
rect 3054 31726 3106 31778
rect 3106 31726 3108 31778
rect 3052 31724 3108 31726
rect 3052 31106 3108 31108
rect 3052 31054 3054 31106
rect 3054 31054 3106 31106
rect 3106 31054 3108 31106
rect 3052 31052 3108 31054
rect 3164 29986 3220 29988
rect 3164 29934 3166 29986
rect 3166 29934 3218 29986
rect 3218 29934 3220 29986
rect 3164 29932 3220 29934
rect 3500 31890 3556 31892
rect 3500 31838 3502 31890
rect 3502 31838 3554 31890
rect 3554 31838 3556 31890
rect 3500 31836 3556 31838
rect 3388 31052 3444 31108
rect 3836 33122 3892 33124
rect 3836 33070 3838 33122
rect 3838 33070 3890 33122
rect 3890 33070 3892 33122
rect 3836 33068 3892 33070
rect 4284 36258 4340 36260
rect 4284 36206 4286 36258
rect 4286 36206 4338 36258
rect 4338 36206 4340 36258
rect 4284 36204 4340 36206
rect 4844 36258 4900 36260
rect 4844 36206 4846 36258
rect 4846 36206 4898 36258
rect 4898 36206 4900 36258
rect 4844 36204 4900 36206
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4396 34300 4452 34356
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4620 33516 4676 33572
rect 5068 33346 5124 33348
rect 5068 33294 5070 33346
rect 5070 33294 5122 33346
rect 5122 33294 5124 33346
rect 5068 33292 5124 33294
rect 3724 30156 3780 30212
rect 2492 27746 2548 27748
rect 2492 27694 2494 27746
rect 2494 27694 2546 27746
rect 2546 27694 2548 27746
rect 2492 27692 2548 27694
rect 2492 25394 2548 25396
rect 2492 25342 2494 25394
rect 2494 25342 2546 25394
rect 2546 25342 2548 25394
rect 2492 25340 2548 25342
rect 2492 23548 2548 23604
rect 2492 21756 2548 21812
rect 3276 29484 3332 29540
rect 3388 29484 3444 29540
rect 5404 34972 5460 35028
rect 5292 34636 5348 34692
rect 5404 34354 5460 34356
rect 5404 34302 5406 34354
rect 5406 34302 5458 34354
rect 5458 34302 5460 34354
rect 5404 34300 5460 34302
rect 4956 32562 5012 32564
rect 4956 32510 4958 32562
rect 4958 32510 5010 32562
rect 5010 32510 5012 32562
rect 4956 32508 5012 32510
rect 3948 31554 4004 31556
rect 3948 31502 3950 31554
rect 3950 31502 4002 31554
rect 4002 31502 4004 31554
rect 3948 31500 4004 31502
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 6412 38668 6468 38724
rect 5628 37772 5684 37828
rect 5964 36370 6020 36372
rect 5964 36318 5966 36370
rect 5966 36318 6018 36370
rect 6018 36318 6020 36370
rect 5964 36316 6020 36318
rect 5628 31948 5684 32004
rect 5964 33346 6020 33348
rect 5964 33294 5966 33346
rect 5966 33294 6018 33346
rect 6018 33294 6020 33346
rect 5964 33292 6020 33294
rect 5964 31836 6020 31892
rect 6300 35084 6356 35140
rect 6188 34914 6244 34916
rect 6188 34862 6190 34914
rect 6190 34862 6242 34914
rect 6242 34862 6244 34914
rect 6188 34860 6244 34862
rect 6972 42028 7028 42084
rect 6972 40460 7028 40516
rect 7420 43650 7476 43652
rect 7420 43598 7422 43650
rect 7422 43598 7474 43650
rect 7474 43598 7476 43650
rect 7420 43596 7476 43598
rect 7308 42140 7364 42196
rect 7084 38946 7140 38948
rect 7084 38894 7086 38946
rect 7086 38894 7138 38946
rect 7138 38894 7140 38946
rect 7084 38892 7140 38894
rect 6748 36370 6804 36372
rect 6748 36318 6750 36370
rect 6750 36318 6802 36370
rect 6802 36318 6804 36370
rect 6748 36316 6804 36318
rect 6412 34188 6468 34244
rect 6748 35196 6804 35252
rect 5516 31500 5572 31556
rect 6524 32284 6580 32340
rect 4396 31106 4452 31108
rect 4396 31054 4398 31106
rect 4398 31054 4450 31106
rect 4450 31054 4452 31106
rect 4396 31052 4452 31054
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4172 30098 4228 30100
rect 4172 30046 4174 30098
rect 4174 30046 4226 30098
rect 4226 30046 4228 30098
rect 4172 30044 4228 30046
rect 5068 30098 5124 30100
rect 5068 30046 5070 30098
rect 5070 30046 5122 30098
rect 5122 30046 5124 30098
rect 5068 30044 5124 30046
rect 4620 29426 4676 29428
rect 4620 29374 4622 29426
rect 4622 29374 4674 29426
rect 4674 29374 4676 29426
rect 4620 29372 4676 29374
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 3388 28588 3444 28644
rect 3948 28642 4004 28644
rect 3948 28590 3950 28642
rect 3950 28590 4002 28642
rect 4002 28590 4004 28642
rect 3948 28588 4004 28590
rect 3276 28530 3332 28532
rect 3276 28478 3278 28530
rect 3278 28478 3330 28530
rect 3330 28478 3332 28530
rect 3276 28476 3332 28478
rect 5852 29986 5908 29988
rect 5852 29934 5854 29986
rect 5854 29934 5906 29986
rect 5906 29934 5908 29986
rect 5852 29932 5908 29934
rect 5740 29820 5796 29876
rect 6076 31276 6132 31332
rect 6188 30268 6244 30324
rect 5740 28588 5796 28644
rect 2940 28364 2996 28420
rect 3500 28418 3556 28420
rect 3500 28366 3502 28418
rect 3502 28366 3554 28418
rect 3554 28366 3556 28418
rect 3500 28364 3556 28366
rect 4732 28252 4788 28308
rect 4172 27970 4228 27972
rect 4172 27918 4174 27970
rect 4174 27918 4226 27970
rect 4226 27918 4228 27970
rect 4172 27916 4228 27918
rect 4956 27970 5012 27972
rect 4956 27918 4958 27970
rect 4958 27918 5010 27970
rect 5010 27918 5012 27970
rect 4956 27916 5012 27918
rect 3724 27244 3780 27300
rect 3500 26796 3556 26852
rect 3724 26850 3780 26852
rect 3724 26798 3726 26850
rect 3726 26798 3778 26850
rect 3778 26798 3780 26850
rect 3724 26796 3780 26798
rect 1708 19964 1764 20020
rect 1708 18172 1764 18228
rect 2492 19964 2548 20020
rect 2492 18172 2548 18228
rect 1708 16380 1764 16436
rect 1820 15708 1876 15764
rect 1708 14588 1764 14644
rect 1708 12850 1764 12852
rect 1708 12798 1710 12850
rect 1710 12798 1762 12850
rect 1762 12798 1764 12850
rect 1708 12796 1764 12798
rect 2492 16380 2548 16436
rect 2492 14588 2548 14644
rect 2044 13356 2100 13412
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 5068 27468 5124 27524
rect 5180 28476 5236 28532
rect 5740 28252 5796 28308
rect 4684 27412 4740 27414
rect 4620 27244 4676 27300
rect 3948 27074 4004 27076
rect 3948 27022 3950 27074
rect 3950 27022 4002 27074
rect 4002 27022 4004 27074
rect 3948 27020 4004 27022
rect 5516 28028 5572 28084
rect 5292 27804 5348 27860
rect 5628 27916 5684 27972
rect 5180 27020 5236 27076
rect 5068 26012 5124 26068
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3836 13356 3892 13412
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2492 12850 2548 12852
rect 2492 12798 2494 12850
rect 2494 12798 2546 12850
rect 2546 12798 2548 12850
rect 2492 12796 2548 12798
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 1708 11004 1764 11060
rect 2492 11004 2548 11060
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2044 9714 2100 9716
rect 2044 9662 2046 9714
rect 2046 9662 2098 9714
rect 2098 9662 2100 9714
rect 2044 9660 2100 9662
rect 1708 9212 1764 9268
rect 2044 9436 2100 9492
rect 2492 9212 2548 9268
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 1708 7980 1764 8036
rect 2492 8034 2548 8036
rect 2492 7982 2494 8034
rect 2494 7982 2546 8034
rect 2546 7982 2548 8034
rect 2492 7980 2548 7982
rect 1708 7420 1764 7476
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 2380 6748 2436 6804
rect 2156 5852 2212 5908
rect 1708 5628 1764 5684
rect 1708 3836 1764 3892
rect 6076 29484 6132 29540
rect 5964 26460 6020 26516
rect 5852 26348 5908 26404
rect 6188 29372 6244 29428
rect 6412 30210 6468 30212
rect 6412 30158 6414 30210
rect 6414 30158 6466 30210
rect 6466 30158 6468 30210
rect 6412 30156 6468 30158
rect 6636 29986 6692 29988
rect 6636 29934 6638 29986
rect 6638 29934 6690 29986
rect 6690 29934 6692 29986
rect 6636 29932 6692 29934
rect 7084 37772 7140 37828
rect 7980 49698 8036 49700
rect 7980 49646 7982 49698
rect 7982 49646 8034 49698
rect 8034 49646 8036 49698
rect 7980 49644 8036 49646
rect 11788 55186 11844 55188
rect 11788 55134 11790 55186
rect 11790 55134 11842 55186
rect 11842 55134 11844 55186
rect 11788 55132 11844 55134
rect 13580 55298 13636 55300
rect 13580 55246 13582 55298
rect 13582 55246 13634 55298
rect 13634 55246 13636 55298
rect 13580 55244 13636 55246
rect 12348 54572 12404 54628
rect 12796 53564 12852 53620
rect 9884 52892 9940 52948
rect 10892 53452 10948 53508
rect 10668 53058 10724 53060
rect 10668 53006 10670 53058
rect 10670 53006 10722 53058
rect 10722 53006 10724 53058
rect 10668 53004 10724 53006
rect 10556 52946 10612 52948
rect 10556 52894 10558 52946
rect 10558 52894 10610 52946
rect 10610 52894 10612 52946
rect 10556 52892 10612 52894
rect 10220 52332 10276 52388
rect 10444 52668 10500 52724
rect 10332 52220 10388 52276
rect 10108 51938 10164 51940
rect 10108 51886 10110 51938
rect 10110 51886 10162 51938
rect 10162 51886 10164 51938
rect 10108 51884 10164 51886
rect 11564 53506 11620 53508
rect 11564 53454 11566 53506
rect 11566 53454 11618 53506
rect 11618 53454 11620 53506
rect 11564 53452 11620 53454
rect 11116 52892 11172 52948
rect 11004 52722 11060 52724
rect 11004 52670 11006 52722
rect 11006 52670 11058 52722
rect 11058 52670 11060 52722
rect 11004 52668 11060 52670
rect 10780 51548 10836 51604
rect 10892 51660 10948 51716
rect 8988 51324 9044 51380
rect 11340 52162 11396 52164
rect 11340 52110 11342 52162
rect 11342 52110 11394 52162
rect 11394 52110 11396 52162
rect 11340 52108 11396 52110
rect 13804 53564 13860 53620
rect 12908 53116 12964 53172
rect 11676 52668 11732 52724
rect 12796 52668 12852 52724
rect 12460 52332 12516 52388
rect 11564 51548 11620 51604
rect 11116 49980 11172 50036
rect 10780 49868 10836 49924
rect 8540 49756 8596 49812
rect 10444 49810 10500 49812
rect 10444 49758 10446 49810
rect 10446 49758 10498 49810
rect 10498 49758 10500 49810
rect 10444 49756 10500 49758
rect 12012 51602 12068 51604
rect 12012 51550 12014 51602
rect 12014 51550 12066 51602
rect 12066 51550 12068 51602
rect 12012 51548 12068 51550
rect 11900 51212 11956 51268
rect 12348 52162 12404 52164
rect 12348 52110 12350 52162
rect 12350 52110 12402 52162
rect 12402 52110 12404 52162
rect 12348 52108 12404 52110
rect 12012 50034 12068 50036
rect 12012 49982 12014 50034
rect 12014 49982 12066 50034
rect 12066 49982 12068 50034
rect 12012 49980 12068 49982
rect 8876 49644 8932 49700
rect 8204 48860 8260 48916
rect 8316 48412 8372 48468
rect 7868 47458 7924 47460
rect 7868 47406 7870 47458
rect 7870 47406 7922 47458
rect 7922 47406 7924 47458
rect 7868 47404 7924 47406
rect 8204 47852 8260 47908
rect 7868 46786 7924 46788
rect 7868 46734 7870 46786
rect 7870 46734 7922 46786
rect 7922 46734 7924 46786
rect 7868 46732 7924 46734
rect 10556 49084 10612 49140
rect 10332 48748 10388 48804
rect 9660 48412 9716 48468
rect 8316 47068 8372 47124
rect 8428 47628 8484 47684
rect 8092 45666 8148 45668
rect 8092 45614 8094 45666
rect 8094 45614 8146 45666
rect 8146 45614 8148 45666
rect 8092 45612 8148 45614
rect 7980 45388 8036 45444
rect 7756 45106 7812 45108
rect 7756 45054 7758 45106
rect 7758 45054 7810 45106
rect 7810 45054 7812 45106
rect 7756 45052 7812 45054
rect 8092 44210 8148 44212
rect 8092 44158 8094 44210
rect 8094 44158 8146 44210
rect 8146 44158 8148 44210
rect 8092 44156 8148 44158
rect 7644 43484 7700 43540
rect 7868 43426 7924 43428
rect 7868 43374 7870 43426
rect 7870 43374 7922 43426
rect 7922 43374 7924 43426
rect 7868 43372 7924 43374
rect 7644 42476 7700 42532
rect 7644 42028 7700 42084
rect 7420 40124 7476 40180
rect 7532 41692 7588 41748
rect 7532 39116 7588 39172
rect 7644 38892 7700 38948
rect 8092 41132 8148 41188
rect 7420 37436 7476 37492
rect 7980 38722 8036 38724
rect 7980 38670 7982 38722
rect 7982 38670 8034 38722
rect 8034 38670 8036 38722
rect 7980 38668 8036 38670
rect 7980 35980 8036 36036
rect 8764 47570 8820 47572
rect 8764 47518 8766 47570
rect 8766 47518 8818 47570
rect 8818 47518 8820 47570
rect 8764 47516 8820 47518
rect 9324 46844 9380 46900
rect 9100 46732 9156 46788
rect 8652 45890 8708 45892
rect 8652 45838 8654 45890
rect 8654 45838 8706 45890
rect 8706 45838 8708 45890
rect 8652 45836 8708 45838
rect 9324 45778 9380 45780
rect 9324 45726 9326 45778
rect 9326 45726 9378 45778
rect 9378 45726 9380 45778
rect 9324 45724 9380 45726
rect 8428 44940 8484 44996
rect 8316 43538 8372 43540
rect 8316 43486 8318 43538
rect 8318 43486 8370 43538
rect 8370 43486 8372 43538
rect 8316 43484 8372 43486
rect 8540 43708 8596 43764
rect 8428 42588 8484 42644
rect 9100 43538 9156 43540
rect 9100 43486 9102 43538
rect 9102 43486 9154 43538
rect 9154 43486 9156 43538
rect 9100 43484 9156 43486
rect 8764 43372 8820 43428
rect 8764 42754 8820 42756
rect 8764 42702 8766 42754
rect 8766 42702 8818 42754
rect 8818 42702 8820 42754
rect 8764 42700 8820 42702
rect 8652 42140 8708 42196
rect 8876 42194 8932 42196
rect 8876 42142 8878 42194
rect 8878 42142 8930 42194
rect 8930 42142 8932 42194
rect 8876 42140 8932 42142
rect 8652 41804 8708 41860
rect 9884 46396 9940 46452
rect 9548 45836 9604 45892
rect 9884 46002 9940 46004
rect 9884 45950 9886 46002
rect 9886 45950 9938 46002
rect 9938 45950 9940 46002
rect 9884 45948 9940 45950
rect 9548 41298 9604 41300
rect 9548 41246 9550 41298
rect 9550 41246 9602 41298
rect 9602 41246 9604 41298
rect 9548 41244 9604 41246
rect 9660 44940 9716 44996
rect 9772 44604 9828 44660
rect 9996 45724 10052 45780
rect 10220 46956 10276 47012
rect 10332 46844 10388 46900
rect 10668 48076 10724 48132
rect 10556 47516 10612 47572
rect 10444 46172 10500 46228
rect 11228 49308 11284 49364
rect 11004 48748 11060 48804
rect 12236 49810 12292 49812
rect 12236 49758 12238 49810
rect 12238 49758 12290 49810
rect 12290 49758 12292 49810
rect 12236 49756 12292 49758
rect 11116 47458 11172 47460
rect 11116 47406 11118 47458
rect 11118 47406 11170 47458
rect 11170 47406 11172 47458
rect 11116 47404 11172 47406
rect 10780 46396 10836 46452
rect 10668 45724 10724 45780
rect 10220 45164 10276 45220
rect 10108 44940 10164 44996
rect 10108 44716 10164 44772
rect 10108 44268 10164 44324
rect 10220 44604 10276 44660
rect 10108 42700 10164 42756
rect 9884 42642 9940 42644
rect 9884 42590 9886 42642
rect 9886 42590 9938 42642
rect 9938 42590 9940 42642
rect 9884 42588 9940 42590
rect 10220 42252 10276 42308
rect 8204 39004 8260 39060
rect 8316 39676 8372 39732
rect 8204 37996 8260 38052
rect 9660 41020 9716 41076
rect 9996 41244 10052 41300
rect 9548 40796 9604 40852
rect 8540 38722 8596 38724
rect 8540 38670 8542 38722
rect 8542 38670 8594 38722
rect 8594 38670 8596 38722
rect 8540 38668 8596 38670
rect 8988 37548 9044 37604
rect 8764 37378 8820 37380
rect 8764 37326 8766 37378
rect 8766 37326 8818 37378
rect 8818 37326 8820 37378
rect 8764 37324 8820 37326
rect 8652 36652 8708 36708
rect 7420 35196 7476 35252
rect 7308 34860 7364 34916
rect 8092 34914 8148 34916
rect 8092 34862 8094 34914
rect 8094 34862 8146 34914
rect 8146 34862 8148 34914
rect 8092 34860 8148 34862
rect 7420 34018 7476 34020
rect 7420 33966 7422 34018
rect 7422 33966 7474 34018
rect 7474 33966 7476 34018
rect 7420 33964 7476 33966
rect 7084 33068 7140 33124
rect 7308 32562 7364 32564
rect 7308 32510 7310 32562
rect 7310 32510 7362 32562
rect 7362 32510 7364 32562
rect 7308 32508 7364 32510
rect 7084 31948 7140 32004
rect 6972 31836 7028 31892
rect 6972 30492 7028 30548
rect 6412 29538 6468 29540
rect 6412 29486 6414 29538
rect 6414 29486 6466 29538
rect 6466 29486 6468 29538
rect 6412 29484 6468 29486
rect 6412 27468 6468 27524
rect 6636 27132 6692 27188
rect 5964 26012 6020 26068
rect 6300 21756 6356 21812
rect 6748 26796 6804 26852
rect 8988 35532 9044 35588
rect 8540 35196 8596 35252
rect 8204 33964 8260 34020
rect 7420 31276 7476 31332
rect 7644 32844 7700 32900
rect 7532 30492 7588 30548
rect 7756 32732 7812 32788
rect 8092 31612 8148 31668
rect 7868 30210 7924 30212
rect 7868 30158 7870 30210
rect 7870 30158 7922 30210
rect 7922 30158 7924 30210
rect 7868 30156 7924 30158
rect 7532 29820 7588 29876
rect 7532 28700 7588 28756
rect 6972 27858 7028 27860
rect 6972 27806 6974 27858
rect 6974 27806 7026 27858
rect 7026 27806 7028 27858
rect 6972 27804 7028 27806
rect 7308 25618 7364 25620
rect 7308 25566 7310 25618
rect 7310 25566 7362 25618
rect 7362 25566 7364 25618
rect 7308 25564 7364 25566
rect 7980 28476 8036 28532
rect 8092 29596 8148 29652
rect 7756 27916 7812 27972
rect 8092 27804 8148 27860
rect 8092 26962 8148 26964
rect 8092 26910 8094 26962
rect 8094 26910 8146 26962
rect 8146 26910 8148 26962
rect 8092 26908 8148 26910
rect 8876 32844 8932 32900
rect 9548 38332 9604 38388
rect 9212 37548 9268 37604
rect 9212 33346 9268 33348
rect 9212 33294 9214 33346
rect 9214 33294 9266 33346
rect 9266 33294 9268 33346
rect 9212 33292 9268 33294
rect 9100 32620 9156 32676
rect 9212 32508 9268 32564
rect 8652 32060 8708 32116
rect 9100 31836 9156 31892
rect 8428 31388 8484 31444
rect 9100 31500 9156 31556
rect 8988 30940 9044 30996
rect 8428 30210 8484 30212
rect 8428 30158 8430 30210
rect 8430 30158 8482 30210
rect 8482 30158 8484 30210
rect 8428 30156 8484 30158
rect 8540 30044 8596 30100
rect 8540 29708 8596 29764
rect 8428 27858 8484 27860
rect 8428 27806 8430 27858
rect 8430 27806 8482 27858
rect 8482 27806 8484 27858
rect 8428 27804 8484 27806
rect 8652 29484 8708 29540
rect 8876 28812 8932 28868
rect 8764 28082 8820 28084
rect 8764 28030 8766 28082
rect 8766 28030 8818 28082
rect 8818 28030 8820 28082
rect 8764 28028 8820 28030
rect 9548 37324 9604 37380
rect 9772 40514 9828 40516
rect 9772 40462 9774 40514
rect 9774 40462 9826 40514
rect 9826 40462 9828 40514
rect 9772 40460 9828 40462
rect 9996 40460 10052 40516
rect 9772 38108 9828 38164
rect 10668 45218 10724 45220
rect 10668 45166 10670 45218
rect 10670 45166 10722 45218
rect 10722 45166 10724 45218
rect 10668 45164 10724 45166
rect 10668 44940 10724 44996
rect 11116 45948 11172 46004
rect 10892 45836 10948 45892
rect 10892 45500 10948 45556
rect 10556 42588 10612 42644
rect 10444 41916 10500 41972
rect 11004 44322 11060 44324
rect 11004 44270 11006 44322
rect 11006 44270 11058 44322
rect 11058 44270 11060 44322
rect 11004 44268 11060 44270
rect 11340 47964 11396 48020
rect 11452 46956 11508 47012
rect 11452 46674 11508 46676
rect 11452 46622 11454 46674
rect 11454 46622 11506 46674
rect 11506 46622 11508 46674
rect 11452 46620 11508 46622
rect 12124 48354 12180 48356
rect 12124 48302 12126 48354
rect 12126 48302 12178 48354
rect 12178 48302 12180 48354
rect 12124 48300 12180 48302
rect 11900 45948 11956 46004
rect 11228 45500 11284 45556
rect 11676 45724 11732 45780
rect 11228 45330 11284 45332
rect 11228 45278 11230 45330
rect 11230 45278 11282 45330
rect 11282 45278 11284 45330
rect 11228 45276 11284 45278
rect 11340 44940 11396 44996
rect 11116 43650 11172 43652
rect 11116 43598 11118 43650
rect 11118 43598 11170 43650
rect 11170 43598 11172 43650
rect 11116 43596 11172 43598
rect 10780 43372 10836 43428
rect 10892 42812 10948 42868
rect 10556 41804 10612 41860
rect 10444 40012 10500 40068
rect 12012 45388 12068 45444
rect 11452 43708 11508 43764
rect 11340 42476 11396 42532
rect 11676 42588 11732 42644
rect 10892 40012 10948 40068
rect 10780 39618 10836 39620
rect 10780 39566 10782 39618
rect 10782 39566 10834 39618
rect 10834 39566 10836 39618
rect 10780 39564 10836 39566
rect 10780 38780 10836 38836
rect 9660 35698 9716 35700
rect 9660 35646 9662 35698
rect 9662 35646 9714 35698
rect 9714 35646 9716 35698
rect 9660 35644 9716 35646
rect 9660 34972 9716 35028
rect 9660 34524 9716 34580
rect 9660 33346 9716 33348
rect 9660 33294 9662 33346
rect 9662 33294 9714 33346
rect 9714 33294 9716 33346
rect 9660 33292 9716 33294
rect 9548 31836 9604 31892
rect 9660 32844 9716 32900
rect 10108 37266 10164 37268
rect 10108 37214 10110 37266
rect 10110 37214 10162 37266
rect 10162 37214 10164 37266
rect 10108 37212 10164 37214
rect 9996 36652 10052 36708
rect 9996 35922 10052 35924
rect 9996 35870 9998 35922
rect 9998 35870 10050 35922
rect 10050 35870 10052 35922
rect 9996 35868 10052 35870
rect 9996 35196 10052 35252
rect 10220 36316 10276 36372
rect 11228 40012 11284 40068
rect 11116 38780 11172 38836
rect 11116 38162 11172 38164
rect 11116 38110 11118 38162
rect 11118 38110 11170 38162
rect 11170 38110 11172 38162
rect 11116 38108 11172 38110
rect 10668 37660 10724 37716
rect 11116 37660 11172 37716
rect 10556 37490 10612 37492
rect 10556 37438 10558 37490
rect 10558 37438 10610 37490
rect 10610 37438 10612 37490
rect 10556 37436 10612 37438
rect 11116 37324 11172 37380
rect 10444 36370 10500 36372
rect 10444 36318 10446 36370
rect 10446 36318 10498 36370
rect 10498 36318 10500 36370
rect 10444 36316 10500 36318
rect 10444 35868 10500 35924
rect 10108 34300 10164 34356
rect 10108 33458 10164 33460
rect 10108 33406 10110 33458
rect 10110 33406 10162 33458
rect 10162 33406 10164 33458
rect 10108 33404 10164 33406
rect 10892 36316 10948 36372
rect 10668 35922 10724 35924
rect 10668 35870 10670 35922
rect 10670 35870 10722 35922
rect 10722 35870 10724 35922
rect 10668 35868 10724 35870
rect 10556 34524 10612 34580
rect 10220 32620 10276 32676
rect 10444 34300 10500 34356
rect 10556 34242 10612 34244
rect 10556 34190 10558 34242
rect 10558 34190 10610 34242
rect 10610 34190 10612 34242
rect 10556 34188 10612 34190
rect 9884 32508 9940 32564
rect 10332 32562 10388 32564
rect 10332 32510 10334 32562
rect 10334 32510 10386 32562
rect 10386 32510 10388 32562
rect 10332 32508 10388 32510
rect 9436 31500 9492 31556
rect 9884 31500 9940 31556
rect 10108 30994 10164 30996
rect 10108 30942 10110 30994
rect 10110 30942 10162 30994
rect 10162 30942 10164 30994
rect 10108 30940 10164 30942
rect 9660 30098 9716 30100
rect 9660 30046 9662 30098
rect 9662 30046 9714 30098
rect 9714 30046 9716 30098
rect 9660 30044 9716 30046
rect 9772 29538 9828 29540
rect 9772 29486 9774 29538
rect 9774 29486 9826 29538
rect 9826 29486 9828 29538
rect 9772 29484 9828 29486
rect 9660 29426 9716 29428
rect 9660 29374 9662 29426
rect 9662 29374 9714 29426
rect 9714 29374 9716 29426
rect 9660 29372 9716 29374
rect 10668 33404 10724 33460
rect 9100 29148 9156 29204
rect 7644 26402 7700 26404
rect 7644 26350 7646 26402
rect 7646 26350 7698 26402
rect 7698 26350 7700 26402
rect 7644 26348 7700 26350
rect 7756 26066 7812 26068
rect 7756 26014 7758 26066
rect 7758 26014 7810 26066
rect 7810 26014 7812 26066
rect 7756 26012 7812 26014
rect 9100 27692 9156 27748
rect 9212 27186 9268 27188
rect 9212 27134 9214 27186
rect 9214 27134 9266 27186
rect 9266 27134 9268 27186
rect 9212 27132 9268 27134
rect 9100 27074 9156 27076
rect 9100 27022 9102 27074
rect 9102 27022 9154 27074
rect 9154 27022 9156 27074
rect 9100 27020 9156 27022
rect 9324 26850 9380 26852
rect 9324 26798 9326 26850
rect 9326 26798 9378 26850
rect 9378 26798 9380 26850
rect 9324 26796 9380 26798
rect 9548 26796 9604 26852
rect 10780 32508 10836 32564
rect 10668 30044 10724 30100
rect 11116 34018 11172 34020
rect 11116 33966 11118 34018
rect 11118 33966 11170 34018
rect 11170 33966 11172 34018
rect 11116 33964 11172 33966
rect 11116 33628 11172 33684
rect 10892 32284 10948 32340
rect 10892 31388 10948 31444
rect 11004 31052 11060 31108
rect 11564 39394 11620 39396
rect 11564 39342 11566 39394
rect 11566 39342 11618 39394
rect 11618 39342 11620 39394
rect 11564 39340 11620 39342
rect 11788 42028 11844 42084
rect 11900 43708 11956 43764
rect 12796 52274 12852 52276
rect 12796 52222 12798 52274
rect 12798 52222 12850 52274
rect 12850 52222 12852 52274
rect 12796 52220 12852 52222
rect 15708 54514 15764 54516
rect 15708 54462 15710 54514
rect 15710 54462 15762 54514
rect 15762 54462 15764 54514
rect 15708 54460 15764 54462
rect 16828 55298 16884 55300
rect 16828 55246 16830 55298
rect 16830 55246 16882 55298
rect 16882 55246 16884 55298
rect 16828 55244 16884 55246
rect 15932 53788 15988 53844
rect 14588 52220 14644 52276
rect 14812 52668 14868 52724
rect 15372 53004 15428 53060
rect 15372 52668 15428 52724
rect 15484 51938 15540 51940
rect 15484 51886 15486 51938
rect 15486 51886 15538 51938
rect 15538 51886 15540 51938
rect 15484 51884 15540 51886
rect 15036 51548 15092 51604
rect 13132 51378 13188 51380
rect 13132 51326 13134 51378
rect 13134 51326 13186 51378
rect 13186 51326 13188 51378
rect 13132 51324 13188 51326
rect 16828 54460 16884 54516
rect 16604 53788 16660 53844
rect 15932 53116 15988 53172
rect 15820 50764 15876 50820
rect 16380 53116 16436 53172
rect 16716 52444 16772 52500
rect 16492 52220 16548 52276
rect 16604 51324 16660 51380
rect 17276 52220 17332 52276
rect 16828 51884 16884 51940
rect 16828 50764 16884 50820
rect 17388 50764 17444 50820
rect 14364 49980 14420 50036
rect 12572 49756 12628 49812
rect 12460 49308 12516 49364
rect 13132 49756 13188 49812
rect 12908 49308 12964 49364
rect 13020 49420 13076 49476
rect 12684 47852 12740 47908
rect 12236 43708 12292 43764
rect 12124 43596 12180 43652
rect 12796 44044 12852 44100
rect 15260 50034 15316 50036
rect 15260 49982 15262 50034
rect 15262 49982 15314 50034
rect 15314 49982 15316 50034
rect 15260 49980 15316 49982
rect 13580 48524 13636 48580
rect 13132 47852 13188 47908
rect 13356 48130 13412 48132
rect 13356 48078 13358 48130
rect 13358 48078 13410 48130
rect 13410 48078 13412 48130
rect 13356 48076 13412 48078
rect 12460 43596 12516 43652
rect 14028 48524 14084 48580
rect 14364 48748 14420 48804
rect 15708 49644 15764 49700
rect 15036 49196 15092 49252
rect 14364 48300 14420 48356
rect 13132 46786 13188 46788
rect 13132 46734 13134 46786
rect 13134 46734 13186 46786
rect 13186 46734 13188 46786
rect 13132 46732 13188 46734
rect 12348 42588 12404 42644
rect 11788 40514 11844 40516
rect 11788 40462 11790 40514
rect 11790 40462 11842 40514
rect 11842 40462 11844 40514
rect 11788 40460 11844 40462
rect 12572 43426 12628 43428
rect 12572 43374 12574 43426
rect 12574 43374 12626 43426
rect 12626 43374 12628 43426
rect 12572 43372 12628 43374
rect 12012 40290 12068 40292
rect 12012 40238 12014 40290
rect 12014 40238 12066 40290
rect 12066 40238 12068 40290
rect 12012 40236 12068 40238
rect 13132 41468 13188 41524
rect 11788 39564 11844 39620
rect 11340 35980 11396 36036
rect 11788 39058 11844 39060
rect 11788 39006 11790 39058
rect 11790 39006 11842 39058
rect 11842 39006 11844 39058
rect 11788 39004 11844 39006
rect 12348 38722 12404 38724
rect 12348 38670 12350 38722
rect 12350 38670 12402 38722
rect 12402 38670 12404 38722
rect 12348 38668 12404 38670
rect 14028 46732 14084 46788
rect 14476 48242 14532 48244
rect 14476 48190 14478 48242
rect 14478 48190 14530 48242
rect 14530 48190 14532 48242
rect 14476 48188 14532 48190
rect 15148 48188 15204 48244
rect 15372 48860 15428 48916
rect 16044 50370 16100 50372
rect 16044 50318 16046 50370
rect 16046 50318 16098 50370
rect 16098 50318 16100 50370
rect 16044 50316 16100 50318
rect 16268 49980 16324 50036
rect 15820 48748 15876 48804
rect 15260 48130 15316 48132
rect 15260 48078 15262 48130
rect 15262 48078 15314 48130
rect 15314 48078 15316 48130
rect 15260 48076 15316 48078
rect 14812 46844 14868 46900
rect 15372 46956 15428 47012
rect 15036 46732 15092 46788
rect 15708 46786 15764 46788
rect 15708 46734 15710 46786
rect 15710 46734 15762 46786
rect 15762 46734 15764 46786
rect 15708 46732 15764 46734
rect 15036 46450 15092 46452
rect 15036 46398 15038 46450
rect 15038 46398 15090 46450
rect 15090 46398 15092 46450
rect 15036 46396 15092 46398
rect 14476 46172 14532 46228
rect 14812 45164 14868 45220
rect 13692 45106 13748 45108
rect 13692 45054 13694 45106
rect 13694 45054 13746 45106
rect 13746 45054 13748 45106
rect 13692 45052 13748 45054
rect 14364 45052 14420 45108
rect 13692 44098 13748 44100
rect 13692 44046 13694 44098
rect 13694 44046 13746 44098
rect 13746 44046 13748 44098
rect 13692 44044 13748 44046
rect 14028 43932 14084 43988
rect 13468 43484 13524 43540
rect 13916 43538 13972 43540
rect 13916 43486 13918 43538
rect 13918 43486 13970 43538
rect 13970 43486 13972 43538
rect 13916 43484 13972 43486
rect 13356 41468 13412 41524
rect 14028 42252 14084 42308
rect 13916 42028 13972 42084
rect 15260 44716 15316 44772
rect 14476 43820 14532 43876
rect 14364 42140 14420 42196
rect 13692 41074 13748 41076
rect 13692 41022 13694 41074
rect 13694 41022 13746 41074
rect 13746 41022 13748 41074
rect 13692 41020 13748 41022
rect 13020 40290 13076 40292
rect 13020 40238 13022 40290
rect 13022 40238 13074 40290
rect 13074 40238 13076 40290
rect 13020 40236 13076 40238
rect 12908 39452 12964 39508
rect 13020 39058 13076 39060
rect 13020 39006 13022 39058
rect 13022 39006 13074 39058
rect 13074 39006 13076 39058
rect 13020 39004 13076 39006
rect 11340 35084 11396 35140
rect 12236 38220 12292 38276
rect 12796 38220 12852 38276
rect 12124 37826 12180 37828
rect 12124 37774 12126 37826
rect 12126 37774 12178 37826
rect 12178 37774 12180 37826
rect 12124 37772 12180 37774
rect 12348 37772 12404 37828
rect 11900 37436 11956 37492
rect 12124 37378 12180 37380
rect 12124 37326 12126 37378
rect 12126 37326 12178 37378
rect 12178 37326 12180 37378
rect 12124 37324 12180 37326
rect 11788 36988 11844 37044
rect 12124 36204 12180 36260
rect 11564 35308 11620 35364
rect 11452 34748 11508 34804
rect 12012 35922 12068 35924
rect 12012 35870 12014 35922
rect 12014 35870 12066 35922
rect 12066 35870 12068 35922
rect 12012 35868 12068 35870
rect 12124 35698 12180 35700
rect 12124 35646 12126 35698
rect 12126 35646 12178 35698
rect 12178 35646 12180 35698
rect 12124 35644 12180 35646
rect 11788 34860 11844 34916
rect 12236 35084 12292 35140
rect 12012 34412 12068 34468
rect 13020 37660 13076 37716
rect 12572 37490 12628 37492
rect 12572 37438 12574 37490
rect 12574 37438 12626 37490
rect 12626 37438 12628 37490
rect 12572 37436 12628 37438
rect 13356 38892 13412 38948
rect 13580 40684 13636 40740
rect 13468 36988 13524 37044
rect 13692 37826 13748 37828
rect 13692 37774 13694 37826
rect 13694 37774 13746 37826
rect 13746 37774 13748 37826
rect 13692 37772 13748 37774
rect 13132 36428 13188 36484
rect 12572 36316 12628 36372
rect 13020 35644 13076 35700
rect 12572 34914 12628 34916
rect 12572 34862 12574 34914
rect 12574 34862 12626 34914
rect 12626 34862 12628 34914
rect 12572 34860 12628 34862
rect 13132 35084 13188 35140
rect 12236 34300 12292 34356
rect 12012 34018 12068 34020
rect 12012 33966 12014 34018
rect 12014 33966 12066 34018
rect 12066 33966 12068 34018
rect 12012 33964 12068 33966
rect 11452 31666 11508 31668
rect 11452 31614 11454 31666
rect 11454 31614 11506 31666
rect 11506 31614 11508 31666
rect 11452 31612 11508 31614
rect 11452 30940 11508 30996
rect 10668 29372 10724 29428
rect 10220 28530 10276 28532
rect 10220 28478 10222 28530
rect 10222 28478 10274 28530
rect 10274 28478 10276 28530
rect 10220 28476 10276 28478
rect 10556 28812 10612 28868
rect 10780 29036 10836 29092
rect 11004 29426 11060 29428
rect 11004 29374 11006 29426
rect 11006 29374 11058 29426
rect 11058 29374 11060 29426
rect 11004 29372 11060 29374
rect 10444 27916 10500 27972
rect 10780 28418 10836 28420
rect 10780 28366 10782 28418
rect 10782 28366 10834 28418
rect 10834 28366 10836 28418
rect 10780 28364 10836 28366
rect 9996 27746 10052 27748
rect 9996 27694 9998 27746
rect 9998 27694 10050 27746
rect 10050 27694 10052 27746
rect 9996 27692 10052 27694
rect 10780 27356 10836 27412
rect 11004 28364 11060 28420
rect 10556 27020 10612 27076
rect 12124 33234 12180 33236
rect 12124 33182 12126 33234
rect 12126 33182 12178 33234
rect 12178 33182 12180 33234
rect 12124 33180 12180 33182
rect 13916 40908 13972 40964
rect 14140 40460 14196 40516
rect 13916 39004 13972 39060
rect 14140 39618 14196 39620
rect 14140 39566 14142 39618
rect 14142 39566 14194 39618
rect 14194 39566 14196 39618
rect 14140 39564 14196 39566
rect 14140 38444 14196 38500
rect 14140 37884 14196 37940
rect 13916 37436 13972 37492
rect 14364 40402 14420 40404
rect 14364 40350 14366 40402
rect 14366 40350 14418 40402
rect 14418 40350 14420 40402
rect 14364 40348 14420 40350
rect 14700 40460 14756 40516
rect 13804 36428 13860 36484
rect 13468 35084 13524 35140
rect 13580 36092 13636 36148
rect 13132 34242 13188 34244
rect 13132 34190 13134 34242
rect 13134 34190 13186 34242
rect 13186 34190 13188 34242
rect 13132 34188 13188 34190
rect 12460 34130 12516 34132
rect 12460 34078 12462 34130
rect 12462 34078 12514 34130
rect 12514 34078 12516 34130
rect 12460 34076 12516 34078
rect 12684 33964 12740 34020
rect 12348 32956 12404 33012
rect 12460 32450 12516 32452
rect 12460 32398 12462 32450
rect 12462 32398 12514 32450
rect 12514 32398 12516 32450
rect 12460 32396 12516 32398
rect 12124 31948 12180 32004
rect 11228 30098 11284 30100
rect 11228 30046 11230 30098
rect 11230 30046 11282 30098
rect 11282 30046 11284 30098
rect 11228 30044 11284 30046
rect 11228 29148 11284 29204
rect 9772 26572 9828 26628
rect 9660 26514 9716 26516
rect 9660 26462 9662 26514
rect 9662 26462 9714 26514
rect 9714 26462 9716 26514
rect 9660 26460 9716 26462
rect 10108 26460 10164 26516
rect 9548 25676 9604 25732
rect 9660 26236 9716 26292
rect 10556 26572 10612 26628
rect 10332 26348 10388 26404
rect 10556 26124 10612 26180
rect 11004 26514 11060 26516
rect 11004 26462 11006 26514
rect 11006 26462 11058 26514
rect 11058 26462 11060 26514
rect 11004 26460 11060 26462
rect 9660 25564 9716 25620
rect 9436 25506 9492 25508
rect 9436 25454 9438 25506
rect 9438 25454 9490 25506
rect 9490 25454 9492 25506
rect 9436 25452 9492 25454
rect 10220 26012 10276 26068
rect 11004 26012 11060 26068
rect 9548 25394 9604 25396
rect 9548 25342 9550 25394
rect 9550 25342 9602 25394
rect 9602 25342 9604 25394
rect 9548 25340 9604 25342
rect 11004 25506 11060 25508
rect 11004 25454 11006 25506
rect 11006 25454 11058 25506
rect 11058 25454 11060 25506
rect 11004 25452 11060 25454
rect 10444 25340 10500 25396
rect 10780 25394 10836 25396
rect 10780 25342 10782 25394
rect 10782 25342 10834 25394
rect 10834 25342 10836 25394
rect 10780 25340 10836 25342
rect 8764 24780 8820 24836
rect 11900 30156 11956 30212
rect 12348 31164 12404 31220
rect 12012 30044 12068 30100
rect 11676 29820 11732 29876
rect 12012 29708 12068 29764
rect 11788 29372 11844 29428
rect 12124 29484 12180 29540
rect 13020 33740 13076 33796
rect 12908 33234 12964 33236
rect 12908 33182 12910 33234
rect 12910 33182 12962 33234
rect 12962 33182 12964 33234
rect 12908 33180 12964 33182
rect 12908 32844 12964 32900
rect 12236 30044 12292 30100
rect 12124 29148 12180 29204
rect 11452 28364 11508 28420
rect 12684 30156 12740 30212
rect 12572 30098 12628 30100
rect 12572 30046 12574 30098
rect 12574 30046 12626 30098
rect 12626 30046 12628 30098
rect 12572 30044 12628 30046
rect 13468 34914 13524 34916
rect 13468 34862 13470 34914
rect 13470 34862 13522 34914
rect 13522 34862 13524 34914
rect 13468 34860 13524 34862
rect 13132 33292 13188 33348
rect 13244 32956 13300 33012
rect 13244 32396 13300 32452
rect 15148 40460 15204 40516
rect 15708 44322 15764 44324
rect 15708 44270 15710 44322
rect 15710 44270 15762 44322
rect 15762 44270 15764 44322
rect 15708 44268 15764 44270
rect 15484 43372 15540 43428
rect 15260 40348 15316 40404
rect 15372 40236 15428 40292
rect 15260 40124 15316 40180
rect 15372 39676 15428 39732
rect 14476 39004 14532 39060
rect 15036 38834 15092 38836
rect 15036 38782 15038 38834
rect 15038 38782 15090 38834
rect 15090 38782 15092 38834
rect 15036 38780 15092 38782
rect 14812 38556 14868 38612
rect 14476 38444 14532 38500
rect 14476 37938 14532 37940
rect 14476 37886 14478 37938
rect 14478 37886 14530 37938
rect 14530 37886 14532 37938
rect 14476 37884 14532 37886
rect 14140 36706 14196 36708
rect 14140 36654 14142 36706
rect 14142 36654 14194 36706
rect 14194 36654 14196 36706
rect 14140 36652 14196 36654
rect 13916 35868 13972 35924
rect 13916 34972 13972 35028
rect 13692 34802 13748 34804
rect 13692 34750 13694 34802
rect 13694 34750 13746 34802
rect 13746 34750 13748 34802
rect 13692 34748 13748 34750
rect 14028 33740 14084 33796
rect 13692 32956 13748 33012
rect 13132 31948 13188 32004
rect 13692 32396 13748 32452
rect 13132 30828 13188 30884
rect 13020 30044 13076 30100
rect 12348 29036 12404 29092
rect 12236 28028 12292 28084
rect 11452 27916 11508 27972
rect 12012 27916 12068 27972
rect 12124 27858 12180 27860
rect 12124 27806 12126 27858
rect 12126 27806 12178 27858
rect 12178 27806 12180 27858
rect 12124 27804 12180 27806
rect 12124 26962 12180 26964
rect 12124 26910 12126 26962
rect 12126 26910 12178 26962
rect 12178 26910 12180 26962
rect 12124 26908 12180 26910
rect 11788 26796 11844 26852
rect 11900 26290 11956 26292
rect 11900 26238 11902 26290
rect 11902 26238 11954 26290
rect 11954 26238 11956 26290
rect 11900 26236 11956 26238
rect 12348 27020 12404 27076
rect 11900 25506 11956 25508
rect 11900 25454 11902 25506
rect 11902 25454 11954 25506
rect 11954 25454 11956 25506
rect 11900 25452 11956 25454
rect 11228 25228 11284 25284
rect 9884 23996 9940 24052
rect 12012 25282 12068 25284
rect 12012 25230 12014 25282
rect 12014 25230 12066 25282
rect 12066 25230 12068 25282
rect 12012 25228 12068 25230
rect 11676 24946 11732 24948
rect 11676 24894 11678 24946
rect 11678 24894 11730 24946
rect 11730 24894 11732 24946
rect 11676 24892 11732 24894
rect 12348 24892 12404 24948
rect 12684 28754 12740 28756
rect 12684 28702 12686 28754
rect 12686 28702 12738 28754
rect 12738 28702 12740 28754
rect 12684 28700 12740 28702
rect 12460 27132 12516 27188
rect 11676 24556 11732 24612
rect 12572 28028 12628 28084
rect 13132 29372 13188 29428
rect 13580 31836 13636 31892
rect 13356 31276 13412 31332
rect 13468 31164 13524 31220
rect 13804 31948 13860 32004
rect 14140 33122 14196 33124
rect 14140 33070 14142 33122
rect 14142 33070 14194 33122
rect 14194 33070 14196 33122
rect 14140 33068 14196 33070
rect 14028 32674 14084 32676
rect 14028 32622 14030 32674
rect 14030 32622 14082 32674
rect 14082 32622 14084 32674
rect 14028 32620 14084 32622
rect 14028 32396 14084 32452
rect 13916 31612 13972 31668
rect 14140 31276 14196 31332
rect 14364 36482 14420 36484
rect 14364 36430 14366 36482
rect 14366 36430 14418 36482
rect 14418 36430 14420 36482
rect 14364 36428 14420 36430
rect 15708 41074 15764 41076
rect 15708 41022 15710 41074
rect 15710 41022 15762 41074
rect 15762 41022 15764 41074
rect 15708 41020 15764 41022
rect 16156 48802 16212 48804
rect 16156 48750 16158 48802
rect 16158 48750 16210 48802
rect 16210 48750 16212 48802
rect 16156 48748 16212 48750
rect 16044 48636 16100 48692
rect 15932 48188 15988 48244
rect 18508 55356 18564 55412
rect 17724 55298 17780 55300
rect 17724 55246 17726 55298
rect 17726 55246 17778 55298
rect 17778 55246 17780 55298
rect 17724 55244 17780 55246
rect 18732 55244 18788 55300
rect 17836 54514 17892 54516
rect 17836 54462 17838 54514
rect 17838 54462 17890 54514
rect 17890 54462 17892 54514
rect 17836 54460 17892 54462
rect 18396 54514 18452 54516
rect 18396 54462 18398 54514
rect 18398 54462 18450 54514
rect 18450 54462 18452 54514
rect 18396 54460 18452 54462
rect 18284 54348 18340 54404
rect 17612 53676 17668 53732
rect 18172 53730 18228 53732
rect 18172 53678 18174 53730
rect 18174 53678 18226 53730
rect 18226 53678 18228 53730
rect 18172 53676 18228 53678
rect 17612 53452 17668 53508
rect 17724 50540 17780 50596
rect 18172 52834 18228 52836
rect 18172 52782 18174 52834
rect 18174 52782 18226 52834
rect 18226 52782 18228 52834
rect 18172 52780 18228 52782
rect 18396 52332 18452 52388
rect 17948 52220 18004 52276
rect 18172 51884 18228 51940
rect 18732 51324 18788 51380
rect 18844 53788 18900 53844
rect 18172 50594 18228 50596
rect 18172 50542 18174 50594
rect 18174 50542 18226 50594
rect 18226 50542 18228 50594
rect 18172 50540 18228 50542
rect 19068 52556 19124 52612
rect 19068 52332 19124 52388
rect 20524 55410 20580 55412
rect 20524 55358 20526 55410
rect 20526 55358 20578 55410
rect 20578 55358 20580 55410
rect 20524 55356 20580 55358
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19964 52780 20020 52836
rect 20748 52220 20804 52276
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 16604 49980 16660 50036
rect 18396 49868 18452 49924
rect 21420 55298 21476 55300
rect 21420 55246 21422 55298
rect 21422 55246 21474 55298
rect 21474 55246 21476 55298
rect 21420 55244 21476 55246
rect 23324 55356 23380 55412
rect 22652 55020 22708 55076
rect 21756 53676 21812 53732
rect 21980 53788 22036 53844
rect 22652 53788 22708 53844
rect 22428 53730 22484 53732
rect 22428 53678 22430 53730
rect 22430 53678 22482 53730
rect 22482 53678 22484 53730
rect 22428 53676 22484 53678
rect 22876 54460 22932 54516
rect 22316 53452 22372 53508
rect 22876 53788 22932 53844
rect 22764 53058 22820 53060
rect 22764 53006 22766 53058
rect 22766 53006 22818 53058
rect 22818 53006 22820 53058
rect 22764 53004 22820 53006
rect 21420 52220 21476 52276
rect 22092 52274 22148 52276
rect 22092 52222 22094 52274
rect 22094 52222 22146 52274
rect 22146 52222 22148 52274
rect 22092 52220 22148 52222
rect 23100 52220 23156 52276
rect 23212 50428 23268 50484
rect 16492 49196 16548 49252
rect 17164 47458 17220 47460
rect 17164 47406 17166 47458
rect 17166 47406 17218 47458
rect 17218 47406 17220 47458
rect 17164 47404 17220 47406
rect 17500 49026 17556 49028
rect 17500 48974 17502 49026
rect 17502 48974 17554 49026
rect 17554 48974 17556 49026
rect 17500 48972 17556 48974
rect 17836 48914 17892 48916
rect 17836 48862 17838 48914
rect 17838 48862 17890 48914
rect 17890 48862 17892 48914
rect 17836 48860 17892 48862
rect 17388 47404 17444 47460
rect 16156 46956 16212 47012
rect 16492 46732 16548 46788
rect 16380 45948 16436 46004
rect 17276 45890 17332 45892
rect 17276 45838 17278 45890
rect 17278 45838 17330 45890
rect 17330 45838 17332 45890
rect 17276 45836 17332 45838
rect 17276 45052 17332 45108
rect 16828 44322 16884 44324
rect 16828 44270 16830 44322
rect 16830 44270 16882 44322
rect 16882 44270 16884 44322
rect 16828 44268 16884 44270
rect 16604 43932 16660 43988
rect 16380 43708 16436 43764
rect 17724 46002 17780 46004
rect 17724 45950 17726 46002
rect 17726 45950 17778 46002
rect 17778 45950 17780 46002
rect 17724 45948 17780 45950
rect 18284 48972 18340 49028
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20524 49196 20580 49252
rect 19068 49026 19124 49028
rect 19068 48974 19070 49026
rect 19070 48974 19122 49026
rect 19122 48974 19124 49026
rect 19068 48972 19124 48974
rect 18508 48524 18564 48580
rect 17948 45724 18004 45780
rect 17612 44434 17668 44436
rect 17612 44382 17614 44434
rect 17614 44382 17666 44434
rect 17666 44382 17668 44434
rect 17612 44380 17668 44382
rect 18172 47292 18228 47348
rect 17500 43762 17556 43764
rect 17500 43710 17502 43762
rect 17502 43710 17554 43762
rect 17554 43710 17556 43762
rect 17500 43708 17556 43710
rect 18060 43708 18116 43764
rect 17612 43650 17668 43652
rect 17612 43598 17614 43650
rect 17614 43598 17666 43650
rect 17666 43598 17668 43650
rect 17612 43596 17668 43598
rect 15932 43484 15988 43540
rect 15036 37660 15092 37716
rect 15036 37212 15092 37268
rect 14924 36652 14980 36708
rect 14812 35810 14868 35812
rect 14812 35758 14814 35810
rect 14814 35758 14866 35810
rect 14866 35758 14868 35810
rect 14812 35756 14868 35758
rect 14700 35196 14756 35252
rect 15148 37042 15204 37044
rect 15148 36990 15150 37042
rect 15150 36990 15202 37042
rect 15202 36990 15204 37042
rect 15148 36988 15204 36990
rect 15596 40348 15652 40404
rect 15708 39452 15764 39508
rect 15820 37826 15876 37828
rect 15820 37774 15822 37826
rect 15822 37774 15874 37826
rect 15874 37774 15876 37826
rect 15820 37772 15876 37774
rect 17724 43372 17780 43428
rect 16716 42194 16772 42196
rect 16716 42142 16718 42194
rect 16718 42142 16770 42194
rect 16770 42142 16772 42194
rect 16716 42140 16772 42142
rect 16604 42082 16660 42084
rect 16604 42030 16606 42082
rect 16606 42030 16658 42082
rect 16658 42030 16660 42082
rect 16604 42028 16660 42030
rect 16380 41132 16436 41188
rect 16156 40684 16212 40740
rect 16492 40236 16548 40292
rect 16380 39452 16436 39508
rect 16492 39340 16548 39396
rect 16044 38108 16100 38164
rect 16156 37884 16212 37940
rect 16156 37548 16212 37604
rect 16492 37548 16548 37604
rect 16044 37324 16100 37380
rect 15932 37266 15988 37268
rect 15932 37214 15934 37266
rect 15934 37214 15986 37266
rect 15986 37214 15988 37266
rect 15932 37212 15988 37214
rect 16492 37378 16548 37380
rect 16492 37326 16494 37378
rect 16494 37326 16546 37378
rect 16546 37326 16548 37378
rect 16492 37324 16548 37326
rect 16156 37212 16212 37268
rect 15484 36764 15540 36820
rect 15260 35756 15316 35812
rect 15148 35532 15204 35588
rect 15372 35586 15428 35588
rect 15372 35534 15374 35586
rect 15374 35534 15426 35586
rect 15426 35534 15428 35586
rect 15372 35532 15428 35534
rect 14364 34412 14420 34468
rect 14364 33068 14420 33124
rect 14364 32674 14420 32676
rect 14364 32622 14366 32674
rect 14366 32622 14418 32674
rect 14418 32622 14420 32674
rect 14364 32620 14420 32622
rect 14924 34802 14980 34804
rect 14924 34750 14926 34802
rect 14926 34750 14978 34802
rect 14978 34750 14980 34802
rect 14924 34748 14980 34750
rect 15148 34748 15204 34804
rect 15036 34524 15092 34580
rect 14700 33964 14756 34020
rect 14812 34412 14868 34468
rect 14588 33122 14644 33124
rect 14588 33070 14590 33122
rect 14590 33070 14642 33122
rect 14642 33070 14644 33122
rect 14588 33068 14644 33070
rect 15260 34412 15316 34468
rect 15260 34130 15316 34132
rect 15260 34078 15262 34130
rect 15262 34078 15314 34130
rect 15314 34078 15316 34130
rect 15260 34076 15316 34078
rect 14924 32732 14980 32788
rect 14252 31164 14308 31220
rect 13804 29820 13860 29876
rect 14028 30044 14084 30100
rect 15036 32284 15092 32340
rect 14924 31948 14980 32004
rect 15148 31948 15204 32004
rect 14812 31666 14868 31668
rect 14812 31614 14814 31666
rect 14814 31614 14866 31666
rect 14866 31614 14868 31666
rect 14812 31612 14868 31614
rect 14924 31554 14980 31556
rect 14924 31502 14926 31554
rect 14926 31502 14978 31554
rect 14978 31502 14980 31554
rect 14924 31500 14980 31502
rect 14700 30716 14756 30772
rect 14812 31276 14868 31332
rect 15148 31218 15204 31220
rect 15148 31166 15150 31218
rect 15150 31166 15202 31218
rect 15202 31166 15204 31218
rect 15148 31164 15204 31166
rect 14812 30604 14868 30660
rect 13692 29538 13748 29540
rect 13692 29486 13694 29538
rect 13694 29486 13746 29538
rect 13746 29486 13748 29538
rect 13692 29484 13748 29486
rect 13356 28700 13412 28756
rect 13916 29372 13972 29428
rect 13692 29036 13748 29092
rect 13132 28028 13188 28084
rect 14140 28140 14196 28196
rect 13692 28028 13748 28084
rect 14028 27692 14084 27748
rect 12796 26684 12852 26740
rect 12796 26514 12852 26516
rect 12796 26462 12798 26514
rect 12798 26462 12850 26514
rect 12850 26462 12852 26514
rect 12796 26460 12852 26462
rect 12572 25394 12628 25396
rect 12572 25342 12574 25394
rect 12574 25342 12626 25394
rect 12626 25342 12628 25394
rect 12572 25340 12628 25342
rect 13580 26962 13636 26964
rect 13580 26910 13582 26962
rect 13582 26910 13634 26962
rect 13634 26910 13636 26962
rect 13580 26908 13636 26910
rect 13244 26514 13300 26516
rect 13244 26462 13246 26514
rect 13246 26462 13298 26514
rect 13298 26462 13300 26514
rect 13244 26460 13300 26462
rect 13692 26514 13748 26516
rect 13692 26462 13694 26514
rect 13694 26462 13746 26514
rect 13746 26462 13748 26514
rect 13692 26460 13748 26462
rect 13580 26236 13636 26292
rect 13020 24892 13076 24948
rect 13132 24668 13188 24724
rect 13356 25116 13412 25172
rect 12460 23772 12516 23828
rect 11340 23548 11396 23604
rect 13692 25282 13748 25284
rect 13692 25230 13694 25282
rect 13694 25230 13746 25282
rect 13746 25230 13748 25282
rect 13692 25228 13748 25230
rect 14364 29820 14420 29876
rect 14924 29708 14980 29764
rect 14812 29596 14868 29652
rect 14364 29426 14420 29428
rect 14364 29374 14366 29426
rect 14366 29374 14418 29426
rect 14418 29374 14420 29426
rect 14364 29372 14420 29374
rect 14476 28924 14532 28980
rect 14812 29372 14868 29428
rect 15484 34188 15540 34244
rect 15820 34076 15876 34132
rect 15484 32450 15540 32452
rect 15484 32398 15486 32450
rect 15486 32398 15538 32450
rect 15538 32398 15540 32450
rect 15484 32396 15540 32398
rect 15708 32396 15764 32452
rect 15484 31724 15540 31780
rect 15484 30828 15540 30884
rect 16156 37042 16212 37044
rect 16156 36990 16158 37042
rect 16158 36990 16210 37042
rect 16210 36990 16212 37042
rect 16156 36988 16212 36990
rect 16380 36988 16436 37044
rect 15932 33852 15988 33908
rect 15932 32956 15988 33012
rect 16828 37772 16884 37828
rect 16604 36988 16660 37044
rect 16828 37436 16884 37492
rect 16604 36316 16660 36372
rect 18396 47458 18452 47460
rect 18396 47406 18398 47458
rect 18398 47406 18450 47458
rect 18450 47406 18452 47458
rect 18396 47404 18452 47406
rect 19964 48972 20020 49028
rect 19628 48914 19684 48916
rect 19628 48862 19630 48914
rect 19630 48862 19682 48914
rect 19682 48862 19684 48914
rect 19628 48860 19684 48862
rect 20412 48914 20468 48916
rect 20412 48862 20414 48914
rect 20414 48862 20466 48914
rect 20466 48862 20468 48914
rect 20412 48860 20468 48862
rect 19740 48748 19796 48804
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19852 48076 19908 48132
rect 19404 47964 19460 48020
rect 19180 47458 19236 47460
rect 19180 47406 19182 47458
rect 19182 47406 19234 47458
rect 19234 47406 19236 47458
rect 19180 47404 19236 47406
rect 18396 44322 18452 44324
rect 18396 44270 18398 44322
rect 18398 44270 18450 44322
rect 18450 44270 18452 44322
rect 18396 44268 18452 44270
rect 18620 44828 18676 44884
rect 18620 43820 18676 43876
rect 18284 43596 18340 43652
rect 18508 43538 18564 43540
rect 18508 43486 18510 43538
rect 18510 43486 18562 43538
rect 18562 43486 18564 43538
rect 18508 43484 18564 43486
rect 17612 42140 17668 42196
rect 17836 42700 17892 42756
rect 18060 42476 18116 42532
rect 18060 42252 18116 42308
rect 17948 42082 18004 42084
rect 17948 42030 17950 42082
rect 17950 42030 18002 42082
rect 18002 42030 18004 42082
rect 17948 42028 18004 42030
rect 18620 42364 18676 42420
rect 18508 42028 18564 42084
rect 17836 41804 17892 41860
rect 17612 41186 17668 41188
rect 17612 41134 17614 41186
rect 17614 41134 17666 41186
rect 17666 41134 17668 41186
rect 17612 41132 17668 41134
rect 17500 40124 17556 40180
rect 17724 40124 17780 40180
rect 17836 40460 17892 40516
rect 17388 39676 17444 39732
rect 17836 39228 17892 39284
rect 18172 40796 18228 40852
rect 18060 40460 18116 40516
rect 18172 39004 18228 39060
rect 18060 38722 18116 38724
rect 18060 38670 18062 38722
rect 18062 38670 18114 38722
rect 18114 38670 18116 38722
rect 18060 38668 18116 38670
rect 19292 46620 19348 46676
rect 20524 48130 20580 48132
rect 20524 48078 20526 48130
rect 20526 48078 20578 48130
rect 20578 48078 20580 48130
rect 20524 48076 20580 48078
rect 20300 47964 20356 48020
rect 20076 47458 20132 47460
rect 20076 47406 20078 47458
rect 20078 47406 20130 47458
rect 20130 47406 20132 47458
rect 20076 47404 20132 47406
rect 20300 47458 20356 47460
rect 20300 47406 20302 47458
rect 20302 47406 20354 47458
rect 20354 47406 20356 47458
rect 20300 47404 20356 47406
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20524 47068 20580 47124
rect 20748 46396 20804 46452
rect 18844 45836 18900 45892
rect 18844 42028 18900 42084
rect 18956 45164 19012 45220
rect 19068 44940 19124 44996
rect 19068 43708 19124 43764
rect 18620 40796 18676 40852
rect 18844 41356 18900 41412
rect 18508 40290 18564 40292
rect 18508 40238 18510 40290
rect 18510 40238 18562 40290
rect 18562 40238 18564 40290
rect 18508 40236 18564 40238
rect 17164 37436 17220 37492
rect 17948 38050 18004 38052
rect 17948 37998 17950 38050
rect 17950 37998 18002 38050
rect 18002 37998 18004 38050
rect 17948 37996 18004 37998
rect 17836 37938 17892 37940
rect 17836 37886 17838 37938
rect 17838 37886 17890 37938
rect 17890 37886 17892 37938
rect 17836 37884 17892 37886
rect 17276 37212 17332 37268
rect 17164 36764 17220 36820
rect 16828 35084 16884 35140
rect 16940 34914 16996 34916
rect 16940 34862 16942 34914
rect 16942 34862 16994 34914
rect 16994 34862 16996 34914
rect 16940 34860 16996 34862
rect 16604 34188 16660 34244
rect 16716 34130 16772 34132
rect 16716 34078 16718 34130
rect 16718 34078 16770 34130
rect 16770 34078 16772 34130
rect 16716 34076 16772 34078
rect 16156 33180 16212 33236
rect 16156 32956 16212 33012
rect 15820 31778 15876 31780
rect 15820 31726 15822 31778
rect 15822 31726 15874 31778
rect 15874 31726 15876 31778
rect 15820 31724 15876 31726
rect 15484 30604 15540 30660
rect 16380 32956 16436 33012
rect 17052 33404 17108 33460
rect 17388 37100 17444 37156
rect 17500 37548 17556 37604
rect 17500 37212 17556 37268
rect 17948 37772 18004 37828
rect 18060 36652 18116 36708
rect 18396 38556 18452 38612
rect 18508 38050 18564 38052
rect 18508 37998 18510 38050
rect 18510 37998 18562 38050
rect 18562 37998 18564 38050
rect 18508 37996 18564 37998
rect 18732 39618 18788 39620
rect 18732 39566 18734 39618
rect 18734 39566 18786 39618
rect 18786 39566 18788 39618
rect 18732 39564 18788 39566
rect 18956 40348 19012 40404
rect 20076 45890 20132 45892
rect 20076 45838 20078 45890
rect 20078 45838 20130 45890
rect 20130 45838 20132 45890
rect 20076 45836 20132 45838
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19516 45164 19572 45220
rect 19964 44716 20020 44772
rect 20748 45388 20804 45444
rect 20860 45948 20916 46004
rect 20748 45164 20804 45220
rect 20524 44994 20580 44996
rect 20524 44942 20526 44994
rect 20526 44942 20578 44994
rect 20578 44942 20580 44994
rect 20524 44940 20580 44942
rect 20300 44156 20356 44212
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19628 43596 19684 43652
rect 20412 42812 20468 42868
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19404 42140 19460 42196
rect 19964 42028 20020 42084
rect 19852 41804 19908 41860
rect 19516 41580 19572 41636
rect 19628 41356 19684 41412
rect 20300 41804 20356 41860
rect 19852 40962 19908 40964
rect 19852 40910 19854 40962
rect 19854 40910 19906 40962
rect 19906 40910 19908 40962
rect 19852 40908 19908 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19292 40402 19348 40404
rect 19292 40350 19294 40402
rect 19294 40350 19346 40402
rect 19346 40350 19348 40402
rect 19292 40348 19348 40350
rect 19628 40348 19684 40404
rect 19180 39116 19236 39172
rect 19292 40124 19348 40180
rect 18844 38722 18900 38724
rect 18844 38670 18846 38722
rect 18846 38670 18898 38722
rect 18898 38670 18900 38722
rect 18844 38668 18900 38670
rect 19404 39788 19460 39844
rect 19404 39228 19460 39284
rect 19292 38780 19348 38836
rect 18284 37436 18340 37492
rect 18396 36876 18452 36932
rect 17836 36258 17892 36260
rect 17836 36206 17838 36258
rect 17838 36206 17890 36258
rect 17890 36206 17892 36258
rect 17836 36204 17892 36206
rect 17276 33516 17332 33572
rect 17052 33180 17108 33236
rect 17164 33068 17220 33124
rect 16268 31218 16324 31220
rect 16268 31166 16270 31218
rect 16270 31166 16322 31218
rect 16322 31166 16324 31218
rect 16268 31164 16324 31166
rect 16828 32674 16884 32676
rect 16828 32622 16830 32674
rect 16830 32622 16882 32674
rect 16882 32622 16884 32674
rect 16828 32620 16884 32622
rect 16044 31052 16100 31108
rect 16044 30828 16100 30884
rect 16268 30828 16324 30884
rect 16156 30156 16212 30212
rect 16156 29932 16212 29988
rect 15708 29650 15764 29652
rect 15708 29598 15710 29650
rect 15710 29598 15762 29650
rect 15762 29598 15764 29650
rect 15708 29596 15764 29598
rect 14924 28418 14980 28420
rect 14924 28366 14926 28418
rect 14926 28366 14978 28418
rect 14978 28366 14980 28418
rect 14924 28364 14980 28366
rect 15260 28924 15316 28980
rect 15148 28252 15204 28308
rect 14700 28028 14756 28084
rect 14364 27356 14420 27412
rect 14476 27074 14532 27076
rect 14476 27022 14478 27074
rect 14478 27022 14530 27074
rect 14530 27022 14532 27074
rect 14476 27020 14532 27022
rect 15484 27858 15540 27860
rect 15484 27806 15486 27858
rect 15486 27806 15538 27858
rect 15538 27806 15540 27858
rect 15484 27804 15540 27806
rect 15820 27580 15876 27636
rect 14924 27356 14980 27412
rect 14364 26908 14420 26964
rect 14252 26572 14308 26628
rect 14028 25452 14084 25508
rect 15708 27356 15764 27412
rect 14924 27020 14980 27076
rect 15148 27074 15204 27076
rect 15148 27022 15150 27074
rect 15150 27022 15202 27074
rect 15202 27022 15204 27074
rect 15148 27020 15204 27022
rect 15372 26962 15428 26964
rect 15372 26910 15374 26962
rect 15374 26910 15426 26962
rect 15426 26910 15428 26962
rect 15372 26908 15428 26910
rect 15036 26402 15092 26404
rect 15036 26350 15038 26402
rect 15038 26350 15090 26402
rect 15090 26350 15092 26402
rect 15036 26348 15092 26350
rect 14924 25618 14980 25620
rect 14924 25566 14926 25618
rect 14926 25566 14978 25618
rect 14978 25566 14980 25618
rect 14924 25564 14980 25566
rect 13804 25116 13860 25172
rect 14028 25004 14084 25060
rect 13916 24722 13972 24724
rect 13916 24670 13918 24722
rect 13918 24670 13970 24722
rect 13970 24670 13972 24722
rect 13916 24668 13972 24670
rect 14700 24892 14756 24948
rect 15596 26684 15652 26740
rect 15484 26460 15540 26516
rect 15708 26402 15764 26404
rect 15708 26350 15710 26402
rect 15710 26350 15762 26402
rect 15762 26350 15764 26402
rect 15708 26348 15764 26350
rect 15260 25564 15316 25620
rect 16268 28082 16324 28084
rect 16268 28030 16270 28082
rect 16270 28030 16322 28082
rect 16322 28030 16324 28082
rect 16268 28028 16324 28030
rect 16492 31948 16548 32004
rect 16604 31388 16660 31444
rect 16828 30604 16884 30660
rect 15932 26684 15988 26740
rect 16604 29036 16660 29092
rect 16604 28364 16660 28420
rect 16716 28252 16772 28308
rect 16716 27634 16772 27636
rect 16716 27582 16718 27634
rect 16718 27582 16770 27634
rect 16770 27582 16772 27634
rect 16716 27580 16772 27582
rect 17724 35420 17780 35476
rect 17724 35196 17780 35252
rect 17500 34242 17556 34244
rect 17500 34190 17502 34242
rect 17502 34190 17554 34242
rect 17554 34190 17556 34242
rect 17500 34188 17556 34190
rect 17612 33964 17668 34020
rect 17276 30492 17332 30548
rect 17612 33404 17668 33460
rect 17836 34972 17892 35028
rect 17836 34636 17892 34692
rect 18060 36482 18116 36484
rect 18060 36430 18062 36482
rect 18062 36430 18114 36482
rect 18114 36430 18116 36482
rect 18060 36428 18116 36430
rect 18396 35868 18452 35924
rect 18396 35532 18452 35588
rect 18284 34748 18340 34804
rect 18844 37996 18900 38052
rect 18508 35084 18564 35140
rect 18508 34636 18564 34692
rect 18620 36652 18676 36708
rect 18060 34524 18116 34580
rect 18508 34354 18564 34356
rect 18508 34302 18510 34354
rect 18510 34302 18562 34354
rect 18562 34302 18564 34354
rect 18508 34300 18564 34302
rect 18956 37772 19012 37828
rect 19068 37884 19124 37940
rect 18844 36594 18900 36596
rect 18844 36542 18846 36594
rect 18846 36542 18898 36594
rect 18898 36542 18900 36594
rect 18844 36540 18900 36542
rect 18956 37324 19012 37380
rect 19180 36876 19236 36932
rect 19292 37996 19348 38052
rect 19180 35810 19236 35812
rect 19180 35758 19182 35810
rect 19182 35758 19234 35810
rect 19234 35758 19236 35810
rect 19180 35756 19236 35758
rect 19404 37548 19460 37604
rect 20748 42082 20804 42084
rect 20748 42030 20750 42082
rect 20750 42030 20802 42082
rect 20802 42030 20804 42082
rect 20748 42028 20804 42030
rect 22764 50204 22820 50260
rect 22204 49868 22260 49924
rect 21756 49698 21812 49700
rect 21756 49646 21758 49698
rect 21758 49646 21810 49698
rect 21810 49646 21812 49698
rect 21756 49644 21812 49646
rect 21532 49196 21588 49252
rect 21868 49026 21924 49028
rect 21868 48974 21870 49026
rect 21870 48974 21922 49026
rect 21922 48974 21924 49026
rect 21868 48972 21924 48974
rect 21420 45836 21476 45892
rect 21532 47404 21588 47460
rect 27916 55970 27972 55972
rect 27916 55918 27918 55970
rect 27918 55918 27970 55970
rect 27970 55918 27972 55970
rect 27916 55916 27972 55918
rect 28588 55916 28644 55972
rect 28364 55804 28420 55860
rect 23436 54460 23492 54516
rect 23660 53842 23716 53844
rect 23660 53790 23662 53842
rect 23662 53790 23714 53842
rect 23714 53790 23716 53842
rect 23660 53788 23716 53790
rect 23548 51996 23604 52052
rect 24780 54348 24836 54404
rect 23548 51436 23604 51492
rect 22428 48300 22484 48356
rect 22092 48188 22148 48244
rect 22316 48188 22372 48244
rect 21644 46956 21700 47012
rect 22092 46674 22148 46676
rect 22092 46622 22094 46674
rect 22094 46622 22146 46674
rect 22146 46622 22148 46674
rect 22092 46620 22148 46622
rect 21868 46284 21924 46340
rect 21756 45778 21812 45780
rect 21756 45726 21758 45778
rect 21758 45726 21810 45778
rect 21810 45726 21812 45778
rect 21756 45724 21812 45726
rect 20972 44882 21028 44884
rect 20972 44830 20974 44882
rect 20974 44830 21026 44882
rect 21026 44830 21028 44882
rect 20972 44828 21028 44830
rect 21420 44268 21476 44324
rect 21420 43932 21476 43988
rect 23212 48412 23268 48468
rect 22876 47180 22932 47236
rect 22988 48300 23044 48356
rect 22652 46956 22708 47012
rect 22316 46172 22372 46228
rect 21868 44156 21924 44212
rect 20972 43820 21028 43876
rect 21756 43484 21812 43540
rect 21756 42866 21812 42868
rect 21756 42814 21758 42866
rect 21758 42814 21810 42866
rect 21810 42814 21812 42866
rect 21756 42812 21812 42814
rect 21308 42530 21364 42532
rect 21308 42478 21310 42530
rect 21310 42478 21362 42530
rect 21362 42478 21364 42530
rect 21308 42476 21364 42478
rect 20972 41804 21028 41860
rect 21532 41692 21588 41748
rect 22092 45836 22148 45892
rect 22428 45778 22484 45780
rect 22428 45726 22430 45778
rect 22430 45726 22482 45778
rect 22482 45726 22484 45778
rect 22428 45724 22484 45726
rect 22092 44716 22148 44772
rect 22204 44380 22260 44436
rect 21980 43820 22036 43876
rect 22092 43932 22148 43988
rect 22204 43762 22260 43764
rect 22204 43710 22206 43762
rect 22206 43710 22258 43762
rect 22258 43710 22260 43762
rect 22204 43708 22260 43710
rect 21980 41970 22036 41972
rect 21980 41918 21982 41970
rect 21982 41918 22034 41970
rect 22034 41918 22036 41970
rect 21980 41916 22036 41918
rect 21420 41186 21476 41188
rect 21420 41134 21422 41186
rect 21422 41134 21474 41186
rect 21474 41134 21476 41186
rect 21420 41132 21476 41134
rect 20524 40908 20580 40964
rect 21084 40908 21140 40964
rect 21532 40348 21588 40404
rect 20636 40124 20692 40180
rect 20412 39564 20468 39620
rect 19628 39506 19684 39508
rect 19628 39454 19630 39506
rect 19630 39454 19682 39506
rect 19682 39454 19684 39506
rect 19628 39452 19684 39454
rect 20300 39340 20356 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19740 38556 19796 38612
rect 21308 39618 21364 39620
rect 21308 39566 21310 39618
rect 21310 39566 21362 39618
rect 21362 39566 21364 39618
rect 21308 39564 21364 39566
rect 21084 39004 21140 39060
rect 19740 38108 19796 38164
rect 20300 38556 20356 38612
rect 19964 38050 20020 38052
rect 19964 37998 19966 38050
rect 19966 37998 20018 38050
rect 20018 37998 20020 38050
rect 19964 37996 20020 37998
rect 19740 37938 19796 37940
rect 19740 37886 19742 37938
rect 19742 37886 19794 37938
rect 19794 37886 19796 37938
rect 19740 37884 19796 37886
rect 20188 37884 20244 37940
rect 19628 37772 19684 37828
rect 19404 37100 19460 37156
rect 19404 35980 19460 36036
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 37324 20132 37380
rect 20076 37100 20132 37156
rect 20300 36988 20356 37044
rect 20860 37660 20916 37716
rect 22204 41692 22260 41748
rect 21980 40908 22036 40964
rect 22204 39564 22260 39620
rect 21980 39058 22036 39060
rect 21980 39006 21982 39058
rect 21982 39006 22034 39058
rect 22034 39006 22036 39058
rect 21980 39004 22036 39006
rect 20748 36540 20804 36596
rect 20860 36428 20916 36484
rect 20188 36370 20244 36372
rect 20188 36318 20190 36370
rect 20190 36318 20242 36370
rect 20242 36318 20244 36370
rect 20188 36316 20244 36318
rect 19740 36258 19796 36260
rect 19740 36206 19742 36258
rect 19742 36206 19794 36258
rect 19794 36206 19796 36258
rect 19740 36204 19796 36206
rect 20412 36204 20468 36260
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 18844 34802 18900 34804
rect 18844 34750 18846 34802
rect 18846 34750 18898 34802
rect 18898 34750 18900 34802
rect 18844 34748 18900 34750
rect 19068 34690 19124 34692
rect 19068 34638 19070 34690
rect 19070 34638 19122 34690
rect 19122 34638 19124 34690
rect 19068 34636 19124 34638
rect 18060 34076 18116 34132
rect 17948 33516 18004 33572
rect 17612 32844 17668 32900
rect 17836 32844 17892 32900
rect 17724 32620 17780 32676
rect 17836 32060 17892 32116
rect 18284 32844 18340 32900
rect 17948 32284 18004 32340
rect 17612 31106 17668 31108
rect 17612 31054 17614 31106
rect 17614 31054 17666 31106
rect 17666 31054 17668 31106
rect 17612 31052 17668 31054
rect 17052 30044 17108 30100
rect 18172 31948 18228 32004
rect 18284 31890 18340 31892
rect 18284 31838 18286 31890
rect 18286 31838 18338 31890
rect 18338 31838 18340 31890
rect 18284 31836 18340 31838
rect 18620 33068 18676 33124
rect 18508 31778 18564 31780
rect 18508 31726 18510 31778
rect 18510 31726 18562 31778
rect 18562 31726 18564 31778
rect 18508 31724 18564 31726
rect 18620 32284 18676 32340
rect 17836 31500 17892 31556
rect 18060 31500 18116 31556
rect 17948 31388 18004 31444
rect 17724 30828 17780 30884
rect 17500 29036 17556 29092
rect 17836 30940 17892 30996
rect 17500 28812 17556 28868
rect 16828 27468 16884 27524
rect 17052 28364 17108 28420
rect 16492 26348 16548 26404
rect 16044 26290 16100 26292
rect 16044 26238 16046 26290
rect 16046 26238 16098 26290
rect 16098 26238 16100 26290
rect 16044 26236 16100 26238
rect 16156 26124 16212 26180
rect 15932 26012 15988 26068
rect 15820 25564 15876 25620
rect 16044 25506 16100 25508
rect 16044 25454 16046 25506
rect 16046 25454 16098 25506
rect 16098 25454 16100 25506
rect 16044 25452 16100 25454
rect 15260 25282 15316 25284
rect 15260 25230 15262 25282
rect 15262 25230 15314 25282
rect 15314 25230 15316 25282
rect 15260 25228 15316 25230
rect 15596 24220 15652 24276
rect 15148 24050 15204 24052
rect 15148 23998 15150 24050
rect 15150 23998 15202 24050
rect 15202 23998 15204 24050
rect 15148 23996 15204 23998
rect 13356 23436 13412 23492
rect 15148 23772 15204 23828
rect 15932 23772 15988 23828
rect 8316 23212 8372 23268
rect 15820 23266 15876 23268
rect 15820 23214 15822 23266
rect 15822 23214 15874 23266
rect 15874 23214 15876 23266
rect 15820 23212 15876 23214
rect 16604 26124 16660 26180
rect 16380 25564 16436 25620
rect 16492 24556 16548 24612
rect 16492 23772 16548 23828
rect 17052 27356 17108 27412
rect 17164 28252 17220 28308
rect 16716 25452 16772 25508
rect 16828 25340 16884 25396
rect 16716 24668 16772 24724
rect 16940 26012 16996 26068
rect 16940 24780 16996 24836
rect 17388 27468 17444 27524
rect 17500 27020 17556 27076
rect 17612 26684 17668 26740
rect 19068 34412 19124 34468
rect 19292 34972 19348 35028
rect 19292 33964 19348 34020
rect 19292 33404 19348 33460
rect 18956 33122 19012 33124
rect 18956 33070 18958 33122
rect 18958 33070 19010 33122
rect 19010 33070 19012 33122
rect 18956 33068 19012 33070
rect 18844 32562 18900 32564
rect 18844 32510 18846 32562
rect 18846 32510 18898 32562
rect 18898 32510 18900 32562
rect 18844 32508 18900 32510
rect 19068 32508 19124 32564
rect 18956 31612 19012 31668
rect 18956 31388 19012 31444
rect 19068 31052 19124 31108
rect 18172 30882 18228 30884
rect 18172 30830 18174 30882
rect 18174 30830 18226 30882
rect 18226 30830 18228 30882
rect 18172 30828 18228 30830
rect 17948 30492 18004 30548
rect 18284 30210 18340 30212
rect 18284 30158 18286 30210
rect 18286 30158 18338 30210
rect 18338 30158 18340 30210
rect 18284 30156 18340 30158
rect 18844 30882 18900 30884
rect 18844 30830 18846 30882
rect 18846 30830 18898 30882
rect 18898 30830 18900 30882
rect 18844 30828 18900 30830
rect 18956 30604 19012 30660
rect 18732 30156 18788 30212
rect 18956 29650 19012 29652
rect 18956 29598 18958 29650
rect 18958 29598 19010 29650
rect 19010 29598 19012 29650
rect 18956 29596 19012 29598
rect 18620 29484 18676 29540
rect 18284 28418 18340 28420
rect 18284 28366 18286 28418
rect 18286 28366 18338 28418
rect 18338 28366 18340 28418
rect 18284 28364 18340 28366
rect 18732 29260 18788 29316
rect 18844 28642 18900 28644
rect 18844 28590 18846 28642
rect 18846 28590 18898 28642
rect 18898 28590 18900 28642
rect 18844 28588 18900 28590
rect 18732 28364 18788 28420
rect 18060 27356 18116 27412
rect 17612 26402 17668 26404
rect 17612 26350 17614 26402
rect 17614 26350 17666 26402
rect 17666 26350 17668 26402
rect 17612 26348 17668 26350
rect 17388 26124 17444 26180
rect 17948 27244 18004 27300
rect 18060 27186 18116 27188
rect 18060 27134 18062 27186
rect 18062 27134 18114 27186
rect 18114 27134 18116 27186
rect 18060 27132 18116 27134
rect 18620 27468 18676 27524
rect 18732 27356 18788 27412
rect 18844 27020 18900 27076
rect 18396 26962 18452 26964
rect 18396 26910 18398 26962
rect 18398 26910 18450 26962
rect 18450 26910 18452 26962
rect 18396 26908 18452 26910
rect 19292 30604 19348 30660
rect 19516 34636 19572 34692
rect 19852 35532 19908 35588
rect 19852 34860 19908 34916
rect 20300 35196 20356 35252
rect 20076 34860 20132 34916
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20412 34524 20468 34580
rect 19516 34018 19572 34020
rect 19516 33966 19518 34018
rect 19518 33966 19570 34018
rect 19570 33966 19572 34018
rect 19516 33964 19572 33966
rect 19516 33404 19572 33460
rect 20076 33628 20132 33684
rect 19852 33404 19908 33460
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 32284 19684 32340
rect 19516 32172 19572 32228
rect 19964 31948 20020 32004
rect 20636 35644 20692 35700
rect 20748 35980 20804 36036
rect 20860 35922 20916 35924
rect 20860 35870 20862 35922
rect 20862 35870 20914 35922
rect 20914 35870 20916 35922
rect 20860 35868 20916 35870
rect 21308 36204 21364 36260
rect 20972 35698 21028 35700
rect 20972 35646 20974 35698
rect 20974 35646 21026 35698
rect 21026 35646 21028 35698
rect 20972 35644 21028 35646
rect 20748 35420 20804 35476
rect 21308 35196 21364 35252
rect 20972 34860 21028 34916
rect 21196 34130 21252 34132
rect 21196 34078 21198 34130
rect 21198 34078 21250 34130
rect 21250 34078 21252 34130
rect 21196 34076 21252 34078
rect 20972 33964 21028 34020
rect 20748 33852 20804 33908
rect 20972 33628 21028 33684
rect 20412 32060 20468 32116
rect 20636 32844 20692 32900
rect 20188 31778 20244 31780
rect 20188 31726 20190 31778
rect 20190 31726 20242 31778
rect 20242 31726 20244 31778
rect 20188 31724 20244 31726
rect 20076 31612 20132 31668
rect 20300 31554 20356 31556
rect 20300 31502 20302 31554
rect 20302 31502 20354 31554
rect 20354 31502 20356 31554
rect 20300 31500 20356 31502
rect 19628 31276 19684 31332
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20076 31106 20132 31108
rect 20076 31054 20078 31106
rect 20078 31054 20130 31106
rect 20130 31054 20132 31106
rect 20076 31052 20132 31054
rect 20748 31612 20804 31668
rect 22092 37548 22148 37604
rect 21644 36876 21700 36932
rect 21532 35980 21588 36036
rect 21756 35308 21812 35364
rect 21420 34076 21476 34132
rect 21644 33964 21700 34020
rect 21532 33346 21588 33348
rect 21532 33294 21534 33346
rect 21534 33294 21586 33346
rect 21586 33294 21588 33346
rect 21532 33292 21588 33294
rect 21980 36258 22036 36260
rect 21980 36206 21982 36258
rect 21982 36206 22034 36258
rect 22034 36206 22036 36258
rect 21980 36204 22036 36206
rect 21644 32956 21700 33012
rect 21756 33852 21812 33908
rect 21308 32060 21364 32116
rect 21420 31948 21476 32004
rect 21420 31388 21476 31444
rect 21644 31948 21700 32004
rect 19516 30716 19572 30772
rect 19292 29932 19348 29988
rect 19404 30044 19460 30100
rect 19628 30268 19684 30324
rect 19964 30716 20020 30772
rect 19964 30380 20020 30436
rect 20860 30604 20916 30660
rect 19964 30044 20020 30100
rect 20412 30098 20468 30100
rect 20412 30046 20414 30098
rect 20414 30046 20466 30098
rect 20466 30046 20468 30098
rect 20412 30044 20468 30046
rect 19516 29650 19572 29652
rect 19516 29598 19518 29650
rect 19518 29598 19570 29650
rect 19570 29598 19572 29650
rect 19516 29596 19572 29598
rect 19292 29036 19348 29092
rect 19292 28642 19348 28644
rect 19292 28590 19294 28642
rect 19294 28590 19346 28642
rect 19346 28590 19348 28642
rect 19292 28588 19348 28590
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20860 29820 20916 29876
rect 20044 29764 20100 29766
rect 19740 29596 19796 29652
rect 21420 30716 21476 30772
rect 21196 30156 21252 30212
rect 20076 29650 20132 29652
rect 20076 29598 20078 29650
rect 20078 29598 20130 29650
rect 20130 29598 20132 29650
rect 20076 29596 20132 29598
rect 20188 29426 20244 29428
rect 20188 29374 20190 29426
rect 20190 29374 20242 29426
rect 20242 29374 20244 29426
rect 20188 29372 20244 29374
rect 19964 29260 20020 29316
rect 20076 28754 20132 28756
rect 20076 28702 20078 28754
rect 20078 28702 20130 28754
rect 20130 28702 20132 28754
rect 20076 28700 20132 28702
rect 20748 29260 20804 29316
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19628 27970 19684 27972
rect 19628 27918 19630 27970
rect 19630 27918 19682 27970
rect 19682 27918 19684 27970
rect 19628 27916 19684 27918
rect 20188 28140 20244 28196
rect 19404 27468 19460 27524
rect 20636 27970 20692 27972
rect 20636 27918 20638 27970
rect 20638 27918 20690 27970
rect 20690 27918 20692 27970
rect 20636 27916 20692 27918
rect 19964 27020 20020 27076
rect 17948 26290 18004 26292
rect 17948 26238 17950 26290
rect 17950 26238 18002 26290
rect 18002 26238 18004 26290
rect 17948 26236 18004 26238
rect 19292 26796 19348 26852
rect 18508 26290 18564 26292
rect 18508 26238 18510 26290
rect 18510 26238 18562 26290
rect 18562 26238 18564 26290
rect 18508 26236 18564 26238
rect 17724 25228 17780 25284
rect 17612 25116 17668 25172
rect 17388 25004 17444 25060
rect 18508 25452 18564 25508
rect 17948 25116 18004 25172
rect 17164 24780 17220 24836
rect 17836 24722 17892 24724
rect 17836 24670 17838 24722
rect 17838 24670 17890 24722
rect 17890 24670 17892 24722
rect 17836 24668 17892 24670
rect 16828 24556 16884 24612
rect 18844 25340 18900 25396
rect 18620 25282 18676 25284
rect 18620 25230 18622 25282
rect 18622 25230 18674 25282
rect 18674 25230 18676 25282
rect 18620 25228 18676 25230
rect 19068 25228 19124 25284
rect 20412 26796 20468 26852
rect 19836 26682 19892 26684
rect 19516 26572 19572 26628
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19964 26012 20020 26068
rect 20412 25900 20468 25956
rect 22092 34972 22148 35028
rect 21980 33516 22036 33572
rect 21980 33234 22036 33236
rect 21980 33182 21982 33234
rect 21982 33182 22034 33234
rect 22034 33182 22036 33234
rect 21980 33180 22036 33182
rect 21868 32844 21924 32900
rect 21868 31724 21924 31780
rect 21980 32508 22036 32564
rect 21868 30604 21924 30660
rect 21980 30380 22036 30436
rect 23436 48188 23492 48244
rect 23100 46674 23156 46676
rect 23100 46622 23102 46674
rect 23102 46622 23154 46674
rect 23154 46622 23156 46674
rect 23100 46620 23156 46622
rect 24444 53452 24500 53508
rect 25116 53788 25172 53844
rect 24892 53452 24948 53508
rect 23996 52892 24052 52948
rect 24780 52668 24836 52724
rect 27580 55074 27636 55076
rect 27580 55022 27582 55074
rect 27582 55022 27634 55074
rect 27634 55022 27636 55074
rect 27580 55020 27636 55022
rect 26012 54402 26068 54404
rect 26012 54350 26014 54402
rect 26014 54350 26066 54402
rect 26066 54350 26068 54402
rect 26012 54348 26068 54350
rect 26348 53842 26404 53844
rect 26348 53790 26350 53842
rect 26350 53790 26402 53842
rect 26402 53790 26404 53842
rect 26348 53788 26404 53790
rect 26572 53788 26628 53844
rect 25564 53506 25620 53508
rect 25564 53454 25566 53506
rect 25566 53454 25618 53506
rect 25618 53454 25620 53506
rect 25564 53452 25620 53454
rect 25452 52946 25508 52948
rect 25452 52894 25454 52946
rect 25454 52894 25506 52946
rect 25506 52894 25508 52946
rect 25452 52892 25508 52894
rect 25228 52332 25284 52388
rect 25228 52108 25284 52164
rect 25452 51996 25508 52052
rect 24556 50540 24612 50596
rect 28140 53788 28196 53844
rect 25900 51212 25956 51268
rect 25452 50540 25508 50596
rect 26236 51996 26292 52052
rect 26460 52556 26516 52612
rect 26460 51996 26516 52052
rect 26012 50540 26068 50596
rect 24668 50370 24724 50372
rect 24668 50318 24670 50370
rect 24670 50318 24722 50370
rect 24722 50318 24724 50370
rect 24668 50316 24724 50318
rect 26684 52892 26740 52948
rect 27020 52946 27076 52948
rect 27020 52894 27022 52946
rect 27022 52894 27074 52946
rect 27074 52894 27076 52946
rect 27020 52892 27076 52894
rect 27020 52220 27076 52276
rect 26684 51996 26740 52052
rect 26684 50652 26740 50708
rect 27356 50706 27412 50708
rect 27356 50654 27358 50706
rect 27358 50654 27410 50706
rect 27410 50654 27412 50706
rect 27356 50652 27412 50654
rect 26796 50594 26852 50596
rect 26796 50542 26798 50594
rect 26798 50542 26850 50594
rect 26850 50542 26852 50594
rect 26796 50540 26852 50542
rect 26236 50204 26292 50260
rect 24332 49420 24388 49476
rect 23884 48412 23940 48468
rect 23548 46620 23604 46676
rect 23660 46396 23716 46452
rect 23324 45330 23380 45332
rect 23324 45278 23326 45330
rect 23326 45278 23378 45330
rect 23378 45278 23380 45330
rect 23324 45276 23380 45278
rect 22988 45164 23044 45220
rect 23660 44940 23716 44996
rect 22652 44380 22708 44436
rect 22652 42812 22708 42868
rect 22540 42754 22596 42756
rect 22540 42702 22542 42754
rect 22542 42702 22594 42754
rect 22594 42702 22596 42754
rect 22540 42700 22596 42702
rect 22428 38780 22484 38836
rect 22652 40626 22708 40628
rect 22652 40574 22654 40626
rect 22654 40574 22706 40626
rect 22706 40574 22708 40626
rect 22652 40572 22708 40574
rect 23100 44716 23156 44772
rect 22876 43484 22932 43540
rect 22876 42700 22932 42756
rect 22876 41858 22932 41860
rect 22876 41806 22878 41858
rect 22878 41806 22930 41858
rect 22930 41806 22932 41858
rect 22876 41804 22932 41806
rect 22876 41298 22932 41300
rect 22876 41246 22878 41298
rect 22878 41246 22930 41298
rect 22930 41246 22932 41298
rect 22876 41244 22932 41246
rect 22428 37938 22484 37940
rect 22428 37886 22430 37938
rect 22430 37886 22482 37938
rect 22482 37886 22484 37938
rect 22428 37884 22484 37886
rect 22540 37324 22596 37380
rect 23436 43932 23492 43988
rect 23100 43148 23156 43204
rect 23996 48188 24052 48244
rect 23884 48076 23940 48132
rect 24220 46674 24276 46676
rect 24220 46622 24222 46674
rect 24222 46622 24274 46674
rect 24274 46622 24276 46674
rect 24220 46620 24276 46622
rect 24108 46284 24164 46340
rect 25788 49698 25844 49700
rect 25788 49646 25790 49698
rect 25790 49646 25842 49698
rect 25842 49646 25844 49698
rect 25788 49644 25844 49646
rect 24668 49026 24724 49028
rect 24668 48974 24670 49026
rect 24670 48974 24722 49026
rect 24722 48974 24724 49026
rect 24668 48972 24724 48974
rect 25340 48524 25396 48580
rect 24556 48242 24612 48244
rect 24556 48190 24558 48242
rect 24558 48190 24610 48242
rect 24610 48190 24612 48242
rect 24556 48188 24612 48190
rect 25452 47516 25508 47572
rect 25564 47292 25620 47348
rect 25228 46674 25284 46676
rect 25228 46622 25230 46674
rect 25230 46622 25282 46674
rect 25282 46622 25284 46674
rect 25228 46620 25284 46622
rect 24892 46284 24948 46340
rect 23996 44604 24052 44660
rect 23884 42700 23940 42756
rect 23100 42028 23156 42084
rect 23436 41916 23492 41972
rect 23100 41692 23156 41748
rect 23100 40684 23156 40740
rect 23212 41186 23268 41188
rect 23212 41134 23214 41186
rect 23214 41134 23266 41186
rect 23266 41134 23268 41186
rect 23212 41132 23268 41134
rect 23212 40572 23268 40628
rect 23436 40572 23492 40628
rect 23100 40402 23156 40404
rect 23100 40350 23102 40402
rect 23102 40350 23154 40402
rect 23154 40350 23156 40402
rect 23100 40348 23156 40350
rect 23772 40348 23828 40404
rect 22764 37548 22820 37604
rect 22988 39116 23044 39172
rect 23996 41916 24052 41972
rect 23996 41132 24052 41188
rect 24556 45778 24612 45780
rect 24556 45726 24558 45778
rect 24558 45726 24610 45778
rect 24610 45726 24612 45778
rect 24556 45724 24612 45726
rect 24668 44994 24724 44996
rect 24668 44942 24670 44994
rect 24670 44942 24722 44994
rect 24722 44942 24724 44994
rect 24668 44940 24724 44942
rect 24444 44604 24500 44660
rect 24668 44380 24724 44436
rect 25340 44994 25396 44996
rect 25340 44942 25342 44994
rect 25342 44942 25394 44994
rect 25394 44942 25396 44994
rect 25340 44940 25396 44942
rect 25116 44604 25172 44660
rect 24780 44210 24836 44212
rect 24780 44158 24782 44210
rect 24782 44158 24834 44210
rect 24834 44158 24836 44210
rect 24780 44156 24836 44158
rect 24332 43932 24388 43988
rect 24668 43538 24724 43540
rect 24668 43486 24670 43538
rect 24670 43486 24722 43538
rect 24722 43486 24724 43538
rect 24668 43484 24724 43486
rect 24332 43036 24388 43092
rect 24668 42978 24724 42980
rect 24668 42926 24670 42978
rect 24670 42926 24722 42978
rect 24722 42926 24724 42978
rect 24668 42924 24724 42926
rect 24556 41916 24612 41972
rect 24332 41244 24388 41300
rect 24780 41970 24836 41972
rect 24780 41918 24782 41970
rect 24782 41918 24834 41970
rect 24834 41918 24836 41970
rect 24780 41916 24836 41918
rect 24780 41244 24836 41300
rect 25228 44322 25284 44324
rect 25228 44270 25230 44322
rect 25230 44270 25282 44322
rect 25282 44270 25284 44322
rect 25228 44268 25284 44270
rect 25116 44210 25172 44212
rect 25116 44158 25118 44210
rect 25118 44158 25170 44210
rect 25170 44158 25172 44210
rect 25116 44156 25172 44158
rect 27580 51212 27636 51268
rect 27132 49026 27188 49028
rect 27132 48974 27134 49026
rect 27134 48974 27186 49026
rect 27186 48974 27188 49026
rect 27132 48972 27188 48974
rect 27356 48636 27412 48692
rect 27468 48524 27524 48580
rect 26572 48242 26628 48244
rect 26572 48190 26574 48242
rect 26574 48190 26626 48242
rect 26626 48190 26628 48242
rect 26572 48188 26628 48190
rect 26908 47516 26964 47572
rect 25900 45164 25956 45220
rect 25788 44994 25844 44996
rect 25788 44942 25790 44994
rect 25790 44942 25842 44994
rect 25842 44942 25844 44994
rect 25788 44940 25844 44942
rect 25788 44604 25844 44660
rect 25116 43372 25172 43428
rect 24780 41074 24836 41076
rect 24780 41022 24782 41074
rect 24782 41022 24834 41074
rect 24834 41022 24836 41074
rect 24780 41020 24836 41022
rect 24780 40460 24836 40516
rect 25004 40124 25060 40180
rect 24668 39788 24724 39844
rect 23324 38780 23380 38836
rect 23212 37996 23268 38052
rect 22988 37324 23044 37380
rect 23100 37548 23156 37604
rect 22652 37100 22708 37156
rect 23100 37100 23156 37156
rect 22876 36370 22932 36372
rect 22876 36318 22878 36370
rect 22878 36318 22930 36370
rect 22930 36318 22932 36370
rect 22876 36316 22932 36318
rect 22876 35868 22932 35924
rect 22540 35644 22596 35700
rect 22764 34748 22820 34804
rect 22652 34636 22708 34692
rect 24220 38946 24276 38948
rect 24220 38894 24222 38946
rect 24222 38894 24274 38946
rect 24274 38894 24276 38946
rect 24220 38892 24276 38894
rect 23324 36876 23380 36932
rect 23436 37660 23492 37716
rect 23660 37212 23716 37268
rect 23436 35420 23492 35476
rect 23660 35196 23716 35252
rect 25452 42252 25508 42308
rect 25676 43148 25732 43204
rect 25676 41970 25732 41972
rect 25676 41918 25678 41970
rect 25678 41918 25730 41970
rect 25730 41918 25732 41970
rect 25676 41916 25732 41918
rect 26124 45106 26180 45108
rect 26124 45054 26126 45106
rect 26126 45054 26178 45106
rect 26178 45054 26180 45106
rect 26124 45052 26180 45054
rect 26348 45164 26404 45220
rect 26124 43372 26180 43428
rect 26236 44322 26292 44324
rect 26236 44270 26238 44322
rect 26238 44270 26290 44322
rect 26290 44270 26292 44322
rect 26236 44268 26292 44270
rect 26348 43372 26404 43428
rect 26236 42364 26292 42420
rect 26348 42252 26404 42308
rect 25788 41580 25844 41636
rect 25900 42028 25956 42084
rect 26348 42082 26404 42084
rect 26348 42030 26350 42082
rect 26350 42030 26402 42082
rect 26402 42030 26404 42082
rect 26348 42028 26404 42030
rect 26236 41970 26292 41972
rect 26236 41918 26238 41970
rect 26238 41918 26290 41970
rect 26290 41918 26292 41970
rect 26236 41916 26292 41918
rect 26236 41356 26292 41412
rect 25900 41020 25956 41076
rect 25340 40178 25396 40180
rect 25340 40126 25342 40178
rect 25342 40126 25394 40178
rect 25394 40126 25396 40178
rect 25340 40124 25396 40126
rect 25452 40012 25508 40068
rect 25452 39788 25508 39844
rect 25564 39452 25620 39508
rect 25564 38722 25620 38724
rect 25564 38670 25566 38722
rect 25566 38670 25618 38722
rect 25618 38670 25620 38722
rect 25564 38668 25620 38670
rect 24108 37772 24164 37828
rect 23884 37660 23940 37716
rect 24444 37436 24500 37492
rect 23884 37378 23940 37380
rect 23884 37326 23886 37378
rect 23886 37326 23938 37378
rect 23938 37326 23940 37378
rect 23884 37324 23940 37326
rect 24556 37548 24612 37604
rect 23884 36652 23940 36708
rect 23996 36540 24052 36596
rect 24220 36540 24276 36596
rect 24108 36482 24164 36484
rect 24108 36430 24110 36482
rect 24110 36430 24162 36482
rect 24162 36430 24164 36482
rect 24108 36428 24164 36430
rect 23772 35084 23828 35140
rect 23548 34972 23604 35028
rect 23772 34748 23828 34804
rect 23548 34524 23604 34580
rect 22204 33068 22260 33124
rect 22316 33180 22372 33236
rect 22428 32732 22484 32788
rect 22428 31778 22484 31780
rect 22428 31726 22430 31778
rect 22430 31726 22482 31778
rect 22482 31726 22484 31778
rect 22428 31724 22484 31726
rect 22204 31612 22260 31668
rect 22652 31164 22708 31220
rect 22428 30492 22484 30548
rect 22540 31052 22596 31108
rect 21308 29596 21364 29652
rect 21980 30098 22036 30100
rect 21980 30046 21982 30098
rect 21982 30046 22034 30098
rect 22034 30046 22036 30098
rect 21980 30044 22036 30046
rect 22428 29932 22484 29988
rect 21756 29426 21812 29428
rect 21756 29374 21758 29426
rect 21758 29374 21810 29426
rect 21810 29374 21812 29426
rect 21756 29372 21812 29374
rect 21644 28252 21700 28308
rect 21532 28140 21588 28196
rect 21644 27132 21700 27188
rect 21420 26908 21476 26964
rect 20076 25228 20132 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 18172 23826 18228 23828
rect 18172 23774 18174 23826
rect 18174 23774 18226 23826
rect 18226 23774 18228 23826
rect 18172 23772 18228 23774
rect 19068 23772 19124 23828
rect 16156 22876 16212 22932
rect 17612 22876 17668 22932
rect 19964 24668 20020 24724
rect 19740 24050 19796 24052
rect 19740 23998 19742 24050
rect 19742 23998 19794 24050
rect 19794 23998 19796 24050
rect 19740 23996 19796 23998
rect 20188 23938 20244 23940
rect 20188 23886 20190 23938
rect 20190 23886 20242 23938
rect 20242 23886 20244 23938
rect 20188 23884 20244 23886
rect 21196 26460 21252 26516
rect 20860 26402 20916 26404
rect 20860 26350 20862 26402
rect 20862 26350 20914 26402
rect 20914 26350 20916 26402
rect 20860 26348 20916 26350
rect 20972 24780 21028 24836
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 21084 23884 21140 23940
rect 21980 26850 22036 26852
rect 21980 26798 21982 26850
rect 21982 26798 22034 26850
rect 22034 26798 22036 26850
rect 21980 26796 22036 26798
rect 21532 25282 21588 25284
rect 21532 25230 21534 25282
rect 21534 25230 21586 25282
rect 21586 25230 21588 25282
rect 21532 25228 21588 25230
rect 22204 29426 22260 29428
rect 22204 29374 22206 29426
rect 22206 29374 22258 29426
rect 22258 29374 22260 29426
rect 22204 29372 22260 29374
rect 22652 29596 22708 29652
rect 22652 28588 22708 28644
rect 22204 26796 22260 26852
rect 22204 26124 22260 26180
rect 21532 24780 21588 24836
rect 21980 24108 22036 24164
rect 22316 24108 22372 24164
rect 22876 33122 22932 33124
rect 22876 33070 22878 33122
rect 22878 33070 22930 33122
rect 22930 33070 22932 33122
rect 22876 33068 22932 33070
rect 22876 32508 22932 32564
rect 22876 31778 22932 31780
rect 22876 31726 22878 31778
rect 22878 31726 22930 31778
rect 22930 31726 22932 31778
rect 22876 31724 22932 31726
rect 22876 31052 22932 31108
rect 22876 30492 22932 30548
rect 23212 33458 23268 33460
rect 23212 33406 23214 33458
rect 23214 33406 23266 33458
rect 23266 33406 23268 33458
rect 23212 33404 23268 33406
rect 23324 33346 23380 33348
rect 23324 33294 23326 33346
rect 23326 33294 23378 33346
rect 23378 33294 23380 33346
rect 23324 33292 23380 33294
rect 23548 33180 23604 33236
rect 23100 32956 23156 33012
rect 23212 33068 23268 33124
rect 23660 33068 23716 33124
rect 24444 36540 24500 36596
rect 24332 35308 24388 35364
rect 24332 34748 24388 34804
rect 23996 34130 24052 34132
rect 23996 34078 23998 34130
rect 23998 34078 24050 34130
rect 24050 34078 24052 34130
rect 23996 34076 24052 34078
rect 23212 31948 23268 32004
rect 23660 31724 23716 31780
rect 23212 30268 23268 30324
rect 23772 30940 23828 30996
rect 23100 30156 23156 30212
rect 22988 28082 23044 28084
rect 22988 28030 22990 28082
rect 22990 28030 23042 28082
rect 23042 28030 23044 28082
rect 22988 28028 23044 28030
rect 22876 27132 22932 27188
rect 23548 29932 23604 29988
rect 23436 29650 23492 29652
rect 23436 29598 23438 29650
rect 23438 29598 23490 29650
rect 23490 29598 23492 29650
rect 23436 29596 23492 29598
rect 23996 30156 24052 30212
rect 23772 29708 23828 29764
rect 23884 30044 23940 30100
rect 23772 29484 23828 29540
rect 24220 31388 24276 31444
rect 25452 36428 25508 36484
rect 25340 35756 25396 35812
rect 25340 35084 25396 35140
rect 24668 33740 24724 33796
rect 24780 33516 24836 33572
rect 24668 32786 24724 32788
rect 24668 32734 24670 32786
rect 24670 32734 24722 32786
rect 24722 32734 24724 32786
rect 24668 32732 24724 32734
rect 25452 34300 25508 34356
rect 25340 33628 25396 33684
rect 25228 33404 25284 33460
rect 25116 33234 25172 33236
rect 25116 33182 25118 33234
rect 25118 33182 25170 33234
rect 25170 33182 25172 33234
rect 25116 33180 25172 33182
rect 25452 32732 25508 32788
rect 25340 32562 25396 32564
rect 25340 32510 25342 32562
rect 25342 32510 25394 32562
rect 25394 32510 25396 32562
rect 25340 32508 25396 32510
rect 24668 30380 24724 30436
rect 24332 30268 24388 30324
rect 24220 29708 24276 29764
rect 23548 29260 23604 29316
rect 23212 28700 23268 28756
rect 23324 28642 23380 28644
rect 23324 28590 23326 28642
rect 23326 28590 23378 28642
rect 23378 28590 23380 28642
rect 23324 28588 23380 28590
rect 23436 28530 23492 28532
rect 23436 28478 23438 28530
rect 23438 28478 23490 28530
rect 23490 28478 23492 28530
rect 23436 28476 23492 28478
rect 23772 27186 23828 27188
rect 23772 27134 23774 27186
rect 23774 27134 23826 27186
rect 23826 27134 23828 27186
rect 23772 27132 23828 27134
rect 24332 29148 24388 29204
rect 24556 28754 24612 28756
rect 24556 28702 24558 28754
rect 24558 28702 24610 28754
rect 24610 28702 24612 28754
rect 24556 28700 24612 28702
rect 24332 28364 24388 28420
rect 24220 28028 24276 28084
rect 24220 27132 24276 27188
rect 23212 26178 23268 26180
rect 23212 26126 23214 26178
rect 23214 26126 23266 26178
rect 23266 26126 23268 26178
rect 23212 26124 23268 26126
rect 22764 25340 22820 25396
rect 23100 25788 23156 25844
rect 22652 25228 22708 25284
rect 23212 25116 23268 25172
rect 23660 26012 23716 26068
rect 22540 24108 22596 24164
rect 23324 24780 23380 24836
rect 22428 23436 22484 23492
rect 21308 23266 21364 23268
rect 21308 23214 21310 23266
rect 21310 23214 21362 23266
rect 21362 23214 21364 23266
rect 21308 23212 21364 23214
rect 23436 25676 23492 25732
rect 24220 25788 24276 25844
rect 24444 25676 24500 25732
rect 23548 25394 23604 25396
rect 23548 25342 23550 25394
rect 23550 25342 23602 25394
rect 23602 25342 23604 25394
rect 23548 25340 23604 25342
rect 24444 25116 24500 25172
rect 23772 24892 23828 24948
rect 24220 24834 24276 24836
rect 24220 24782 24222 24834
rect 24222 24782 24274 24834
rect 24274 24782 24276 24834
rect 24220 24780 24276 24782
rect 24444 23996 24500 24052
rect 24668 27746 24724 27748
rect 24668 27694 24670 27746
rect 24670 27694 24722 27746
rect 24722 27694 24724 27746
rect 24668 27692 24724 27694
rect 25004 30210 25060 30212
rect 25004 30158 25006 30210
rect 25006 30158 25058 30210
rect 25058 30158 25060 30210
rect 25004 30156 25060 30158
rect 25116 30940 25172 30996
rect 25564 31948 25620 32004
rect 25116 30268 25172 30324
rect 25228 29932 25284 29988
rect 25116 28642 25172 28644
rect 25116 28590 25118 28642
rect 25118 28590 25170 28642
rect 25170 28590 25172 28642
rect 25116 28588 25172 28590
rect 25228 27074 25284 27076
rect 25228 27022 25230 27074
rect 25230 27022 25282 27074
rect 25282 27022 25284 27074
rect 25228 27020 25284 27022
rect 25228 26572 25284 26628
rect 25788 39788 25844 39844
rect 26124 39788 26180 39844
rect 26348 39452 26404 39508
rect 26236 38946 26292 38948
rect 26236 38894 26238 38946
rect 26238 38894 26290 38946
rect 26290 38894 26292 38946
rect 26236 38892 26292 38894
rect 25788 37548 25844 37604
rect 25788 37378 25844 37380
rect 25788 37326 25790 37378
rect 25790 37326 25842 37378
rect 25842 37326 25844 37378
rect 25788 37324 25844 37326
rect 25788 36988 25844 37044
rect 26124 38050 26180 38052
rect 26124 37998 26126 38050
rect 26126 37998 26178 38050
rect 26178 37998 26180 38050
rect 26124 37996 26180 37998
rect 26124 37436 26180 37492
rect 25900 36540 25956 36596
rect 25788 35420 25844 35476
rect 26012 34748 26068 34804
rect 27916 49026 27972 49028
rect 27916 48974 27918 49026
rect 27918 48974 27970 49026
rect 27970 48974 27972 49026
rect 27916 48972 27972 48974
rect 27692 47404 27748 47460
rect 27804 48636 27860 48692
rect 27580 46956 27636 47012
rect 28252 51266 28308 51268
rect 28252 51214 28254 51266
rect 28254 51214 28306 51266
rect 28306 51214 28308 51266
rect 28252 51212 28308 51214
rect 29260 55298 29316 55300
rect 29260 55246 29262 55298
rect 29262 55246 29314 55298
rect 29314 55246 29316 55298
rect 29260 55244 29316 55246
rect 29148 54626 29204 54628
rect 29148 54574 29150 54626
rect 29150 54574 29202 54626
rect 29202 54574 29204 54626
rect 29148 54572 29204 54574
rect 28812 54514 28868 54516
rect 28812 54462 28814 54514
rect 28814 54462 28866 54514
rect 28866 54462 28868 54514
rect 28812 54460 28868 54462
rect 31836 54626 31892 54628
rect 31836 54574 31838 54626
rect 31838 54574 31890 54626
rect 31890 54574 31892 54626
rect 31836 54572 31892 54574
rect 29260 53900 29316 53956
rect 29148 53452 29204 53508
rect 30044 54514 30100 54516
rect 30044 54462 30046 54514
rect 30046 54462 30098 54514
rect 30098 54462 30100 54514
rect 30044 54460 30100 54462
rect 30380 53788 30436 53844
rect 30156 53452 30212 53508
rect 29932 53058 29988 53060
rect 29932 53006 29934 53058
rect 29934 53006 29986 53058
rect 29986 53006 29988 53058
rect 29932 53004 29988 53006
rect 33180 55244 33236 55300
rect 32508 55020 32564 55076
rect 32508 54572 32564 54628
rect 32060 53676 32116 53732
rect 32620 53618 32676 53620
rect 32620 53566 32622 53618
rect 32622 53566 32674 53618
rect 32674 53566 32676 53618
rect 32620 53564 32676 53566
rect 32172 53058 32228 53060
rect 32172 53006 32174 53058
rect 32174 53006 32226 53058
rect 32226 53006 32228 53058
rect 32172 53004 32228 53006
rect 30716 52946 30772 52948
rect 30716 52894 30718 52946
rect 30718 52894 30770 52946
rect 30770 52894 30772 52946
rect 30716 52892 30772 52894
rect 31836 52892 31892 52948
rect 29372 52162 29428 52164
rect 29372 52110 29374 52162
rect 29374 52110 29426 52162
rect 29426 52110 29428 52162
rect 29372 52108 29428 52110
rect 33404 54626 33460 54628
rect 33404 54574 33406 54626
rect 33406 54574 33458 54626
rect 33458 54574 33460 54626
rect 33404 54572 33460 54574
rect 33628 54572 33684 54628
rect 33068 53564 33124 53620
rect 33292 53788 33348 53844
rect 33180 53116 33236 53172
rect 29484 51996 29540 52052
rect 32732 52274 32788 52276
rect 32732 52222 32734 52274
rect 32734 52222 32786 52274
rect 32786 52222 32788 52274
rect 32732 52220 32788 52222
rect 33852 54460 33908 54516
rect 33628 53788 33684 53844
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 36092 54684 36148 54740
rect 33964 54348 34020 54404
rect 33852 53564 33908 53620
rect 34636 53564 34692 53620
rect 33852 52946 33908 52948
rect 33852 52894 33854 52946
rect 33854 52894 33906 52946
rect 33906 52894 33908 52946
rect 33852 52892 33908 52894
rect 32620 51212 32676 51268
rect 28028 48524 28084 48580
rect 28140 49084 28196 49140
rect 27356 45778 27412 45780
rect 27356 45726 27358 45778
rect 27358 45726 27410 45778
rect 27410 45726 27412 45778
rect 27356 45724 27412 45726
rect 26572 44210 26628 44212
rect 26572 44158 26574 44210
rect 26574 44158 26626 44210
rect 26626 44158 26628 44210
rect 26572 44156 26628 44158
rect 26572 43932 26628 43988
rect 26684 43484 26740 43540
rect 27244 43484 27300 43540
rect 27132 42924 27188 42980
rect 27020 42252 27076 42308
rect 26572 41970 26628 41972
rect 26572 41918 26574 41970
rect 26574 41918 26626 41970
rect 26626 41918 26628 41970
rect 26572 41916 26628 41918
rect 26908 41356 26964 41412
rect 26796 41020 26852 41076
rect 26684 40908 26740 40964
rect 26908 40348 26964 40404
rect 27020 39340 27076 39396
rect 26572 38722 26628 38724
rect 26572 38670 26574 38722
rect 26574 38670 26626 38722
rect 26626 38670 26628 38722
rect 26572 38668 26628 38670
rect 26908 38834 26964 38836
rect 26908 38782 26910 38834
rect 26910 38782 26962 38834
rect 26962 38782 26964 38834
rect 26908 38780 26964 38782
rect 27244 40348 27300 40404
rect 27804 42588 27860 42644
rect 27580 41356 27636 41412
rect 30268 50764 30324 50820
rect 28588 49308 28644 49364
rect 29260 48860 29316 48916
rect 28588 48076 28644 48132
rect 28700 48636 28756 48692
rect 28476 47516 28532 47572
rect 28140 44380 28196 44436
rect 29036 48242 29092 48244
rect 29036 48190 29038 48242
rect 29038 48190 29090 48242
rect 29090 48190 29092 48242
rect 29036 48188 29092 48190
rect 28700 47516 28756 47572
rect 28812 45612 28868 45668
rect 28252 43372 28308 43428
rect 28476 42700 28532 42756
rect 27580 41132 27636 41188
rect 28140 41298 28196 41300
rect 28140 41246 28142 41298
rect 28142 41246 28194 41298
rect 28194 41246 28196 41298
rect 28140 41244 28196 41246
rect 28588 42140 28644 42196
rect 28700 41916 28756 41972
rect 28588 41468 28644 41524
rect 28476 40908 28532 40964
rect 28252 40402 28308 40404
rect 28252 40350 28254 40402
rect 28254 40350 28306 40402
rect 28306 40350 28308 40402
rect 28252 40348 28308 40350
rect 29148 45164 29204 45220
rect 29148 44380 29204 44436
rect 29148 43650 29204 43652
rect 29148 43598 29150 43650
rect 29150 43598 29202 43650
rect 29202 43598 29204 43650
rect 29148 43596 29204 43598
rect 32508 49980 32564 50036
rect 30604 49084 30660 49140
rect 32060 49084 32116 49140
rect 29820 48354 29876 48356
rect 29820 48302 29822 48354
rect 29822 48302 29874 48354
rect 29874 48302 29876 48354
rect 29820 48300 29876 48302
rect 30268 47852 30324 47908
rect 29484 45836 29540 45892
rect 29372 45276 29428 45332
rect 30156 46956 30212 47012
rect 31500 48242 31556 48244
rect 31500 48190 31502 48242
rect 31502 48190 31554 48242
rect 31554 48190 31556 48242
rect 31500 48188 31556 48190
rect 32060 48860 32116 48916
rect 31836 48748 31892 48804
rect 32172 48188 32228 48244
rect 31612 47964 31668 48020
rect 31724 48076 31780 48132
rect 31164 47628 31220 47684
rect 30940 47516 30996 47572
rect 31276 47458 31332 47460
rect 31276 47406 31278 47458
rect 31278 47406 31330 47458
rect 31330 47406 31332 47458
rect 31276 47404 31332 47406
rect 30268 46844 30324 46900
rect 31612 47068 31668 47124
rect 30044 46172 30100 46228
rect 29820 44604 29876 44660
rect 29932 44546 29988 44548
rect 29932 44494 29934 44546
rect 29934 44494 29986 44546
rect 29986 44494 29988 44546
rect 29932 44492 29988 44494
rect 29820 42754 29876 42756
rect 29820 42702 29822 42754
rect 29822 42702 29874 42754
rect 29874 42702 29876 42754
rect 29820 42700 29876 42702
rect 30940 44492 30996 44548
rect 30380 44380 30436 44436
rect 30604 43932 30660 43988
rect 30268 43484 30324 43540
rect 27692 40012 27748 40068
rect 27804 40290 27860 40292
rect 27804 40238 27806 40290
rect 27806 40238 27858 40290
rect 27858 40238 27860 40290
rect 27804 40236 27860 40238
rect 27468 38892 27524 38948
rect 29372 41356 29428 41412
rect 29148 41244 29204 41300
rect 27916 40124 27972 40180
rect 29372 40796 29428 40852
rect 28588 39788 28644 39844
rect 28028 39618 28084 39620
rect 28028 39566 28030 39618
rect 28030 39566 28082 39618
rect 28082 39566 28084 39618
rect 28028 39564 28084 39566
rect 26684 37938 26740 37940
rect 26684 37886 26686 37938
rect 26686 37886 26738 37938
rect 26738 37886 26740 37938
rect 26684 37884 26740 37886
rect 26460 37266 26516 37268
rect 26460 37214 26462 37266
rect 26462 37214 26514 37266
rect 26514 37214 26516 37266
rect 26460 37212 26516 37214
rect 26684 35586 26740 35588
rect 26684 35534 26686 35586
rect 26686 35534 26738 35586
rect 26738 35534 26740 35586
rect 26684 35532 26740 35534
rect 26684 35308 26740 35364
rect 26236 34972 26292 35028
rect 26908 37548 26964 37604
rect 26908 37212 26964 37268
rect 27020 35868 27076 35924
rect 26908 35756 26964 35812
rect 26908 35308 26964 35364
rect 26236 34188 26292 34244
rect 26348 33852 26404 33908
rect 27132 35586 27188 35588
rect 27132 35534 27134 35586
rect 27134 35534 27186 35586
rect 27186 35534 27188 35586
rect 27132 35532 27188 35534
rect 27132 35308 27188 35364
rect 27132 34972 27188 35028
rect 27020 34636 27076 34692
rect 27356 37884 27412 37940
rect 28252 38668 28308 38724
rect 28140 38556 28196 38612
rect 28028 38444 28084 38500
rect 27580 37772 27636 37828
rect 26572 33740 26628 33796
rect 26460 33628 26516 33684
rect 26012 32620 26068 32676
rect 26796 33570 26852 33572
rect 26796 33518 26798 33570
rect 26798 33518 26850 33570
rect 26850 33518 26852 33570
rect 26796 33516 26852 33518
rect 27020 33292 27076 33348
rect 26908 33180 26964 33236
rect 26684 31388 26740 31444
rect 26348 30828 26404 30884
rect 25452 30044 25508 30100
rect 25788 30156 25844 30212
rect 25900 30098 25956 30100
rect 25900 30046 25902 30098
rect 25902 30046 25954 30098
rect 25954 30046 25956 30098
rect 25900 30044 25956 30046
rect 26796 30940 26852 30996
rect 26460 30156 26516 30212
rect 27244 34018 27300 34020
rect 27244 33966 27246 34018
rect 27246 33966 27298 34018
rect 27298 33966 27300 34018
rect 27244 33964 27300 33966
rect 27244 33628 27300 33684
rect 27468 37548 27524 37604
rect 27916 38332 27972 38388
rect 27804 37154 27860 37156
rect 27804 37102 27806 37154
rect 27806 37102 27858 37154
rect 27858 37102 27860 37154
rect 27804 37100 27860 37102
rect 27580 36594 27636 36596
rect 27580 36542 27582 36594
rect 27582 36542 27634 36594
rect 27634 36542 27636 36594
rect 27580 36540 27636 36542
rect 29036 38722 29092 38724
rect 29036 38670 29038 38722
rect 29038 38670 29090 38722
rect 29090 38670 29092 38722
rect 29036 38668 29092 38670
rect 29820 40290 29876 40292
rect 29820 40238 29822 40290
rect 29822 40238 29874 40290
rect 29874 40238 29876 40290
rect 29820 40236 29876 40238
rect 29596 40012 29652 40068
rect 30156 41468 30212 41524
rect 30604 42700 30660 42756
rect 30492 42364 30548 42420
rect 30940 43484 30996 43540
rect 30492 40402 30548 40404
rect 30492 40350 30494 40402
rect 30494 40350 30546 40402
rect 30546 40350 30548 40402
rect 30492 40348 30548 40350
rect 30268 39842 30324 39844
rect 30268 39790 30270 39842
rect 30270 39790 30322 39842
rect 30322 39790 30324 39842
rect 30268 39788 30324 39790
rect 28588 38220 28644 38276
rect 29260 38332 29316 38388
rect 28140 37884 28196 37940
rect 28476 37548 28532 37604
rect 28028 36316 28084 36372
rect 27580 35756 27636 35812
rect 27804 35698 27860 35700
rect 27804 35646 27806 35698
rect 27806 35646 27858 35698
rect 27858 35646 27860 35698
rect 27804 35644 27860 35646
rect 27804 35308 27860 35364
rect 28028 35308 28084 35364
rect 28476 37100 28532 37156
rect 28700 37884 28756 37940
rect 29708 37826 29764 37828
rect 29708 37774 29710 37826
rect 29710 37774 29762 37826
rect 29762 37774 29764 37826
rect 29708 37772 29764 37774
rect 29036 37490 29092 37492
rect 29036 37438 29038 37490
rect 29038 37438 29090 37490
rect 29090 37438 29092 37490
rect 29036 37436 29092 37438
rect 29484 37490 29540 37492
rect 29484 37438 29486 37490
rect 29486 37438 29538 37490
rect 29538 37438 29540 37490
rect 29484 37436 29540 37438
rect 29596 37378 29652 37380
rect 29596 37326 29598 37378
rect 29598 37326 29650 37378
rect 29650 37326 29652 37378
rect 29596 37324 29652 37326
rect 28924 37212 28980 37268
rect 28364 36370 28420 36372
rect 28364 36318 28366 36370
rect 28366 36318 28418 36370
rect 28418 36318 28420 36370
rect 28364 36316 28420 36318
rect 28476 36258 28532 36260
rect 28476 36206 28478 36258
rect 28478 36206 28530 36258
rect 28530 36206 28532 36258
rect 28476 36204 28532 36206
rect 28700 35922 28756 35924
rect 28700 35870 28702 35922
rect 28702 35870 28754 35922
rect 28754 35870 28756 35922
rect 28700 35868 28756 35870
rect 28252 35698 28308 35700
rect 28252 35646 28254 35698
rect 28254 35646 28306 35698
rect 28306 35646 28308 35698
rect 28252 35644 28308 35646
rect 28140 35084 28196 35140
rect 28252 34914 28308 34916
rect 28252 34862 28254 34914
rect 28254 34862 28306 34914
rect 28306 34862 28308 34914
rect 28252 34860 28308 34862
rect 27692 34690 27748 34692
rect 27692 34638 27694 34690
rect 27694 34638 27746 34690
rect 27746 34638 27748 34690
rect 27692 34636 27748 34638
rect 28140 34636 28196 34692
rect 29820 37266 29876 37268
rect 29820 37214 29822 37266
rect 29822 37214 29874 37266
rect 29874 37214 29876 37266
rect 29820 37212 29876 37214
rect 29596 37100 29652 37156
rect 29148 36652 29204 36708
rect 29260 36258 29316 36260
rect 29260 36206 29262 36258
rect 29262 36206 29314 36258
rect 29314 36206 29316 36258
rect 29260 36204 29316 36206
rect 29148 35308 29204 35364
rect 29036 35084 29092 35140
rect 28028 34242 28084 34244
rect 28028 34190 28030 34242
rect 28030 34190 28082 34242
rect 28082 34190 28084 34242
rect 28028 34188 28084 34190
rect 27580 33906 27636 33908
rect 27580 33854 27582 33906
rect 27582 33854 27634 33906
rect 27634 33854 27636 33906
rect 27580 33852 27636 33854
rect 27244 33180 27300 33236
rect 27468 32844 27524 32900
rect 27692 33516 27748 33572
rect 27804 33964 27860 34020
rect 28252 34524 28308 34580
rect 28252 33964 28308 34020
rect 28700 33852 28756 33908
rect 28476 33516 28532 33572
rect 28028 33346 28084 33348
rect 28028 33294 28030 33346
rect 28030 33294 28082 33346
rect 28082 33294 28084 33346
rect 28028 33292 28084 33294
rect 28252 33234 28308 33236
rect 28252 33182 28254 33234
rect 28254 33182 28306 33234
rect 28306 33182 28308 33234
rect 28252 33180 28308 33182
rect 27580 32620 27636 32676
rect 27692 33122 27748 33124
rect 27692 33070 27694 33122
rect 27694 33070 27746 33122
rect 27746 33070 27748 33122
rect 27692 33068 27748 33070
rect 28812 33292 28868 33348
rect 28364 32674 28420 32676
rect 28364 32622 28366 32674
rect 28366 32622 28418 32674
rect 28418 32622 28420 32674
rect 28364 32620 28420 32622
rect 27692 32284 27748 32340
rect 27132 31276 27188 31332
rect 25452 28364 25508 28420
rect 26348 29036 26404 29092
rect 26236 28924 26292 28980
rect 26684 28812 26740 28868
rect 26908 28924 26964 28980
rect 26012 28642 26068 28644
rect 26012 28590 26014 28642
rect 26014 28590 26066 28642
rect 26066 28590 26068 28642
rect 26012 28588 26068 28590
rect 25676 27692 25732 27748
rect 25900 27580 25956 27636
rect 25900 27020 25956 27076
rect 26460 27858 26516 27860
rect 26460 27806 26462 27858
rect 26462 27806 26514 27858
rect 26514 27806 26516 27858
rect 26460 27804 26516 27806
rect 26684 27916 26740 27972
rect 28028 31666 28084 31668
rect 28028 31614 28030 31666
rect 28030 31614 28082 31666
rect 28082 31614 28084 31666
rect 28028 31612 28084 31614
rect 28476 31388 28532 31444
rect 29260 34690 29316 34692
rect 29260 34638 29262 34690
rect 29262 34638 29314 34690
rect 29314 34638 29316 34690
rect 29260 34636 29316 34638
rect 29372 34188 29428 34244
rect 29260 34018 29316 34020
rect 29260 33966 29262 34018
rect 29262 33966 29314 34018
rect 29314 33966 29316 34018
rect 29260 33964 29316 33966
rect 29484 33964 29540 34020
rect 29260 33234 29316 33236
rect 29260 33182 29262 33234
rect 29262 33182 29314 33234
rect 29314 33182 29316 33234
rect 29260 33180 29316 33182
rect 29148 33068 29204 33124
rect 27692 30994 27748 30996
rect 27692 30942 27694 30994
rect 27694 30942 27746 30994
rect 27746 30942 27748 30994
rect 27692 30940 27748 30942
rect 27916 30716 27972 30772
rect 28028 30156 28084 30212
rect 27244 29650 27300 29652
rect 27244 29598 27246 29650
rect 27246 29598 27298 29650
rect 27298 29598 27300 29650
rect 27244 29596 27300 29598
rect 27804 29650 27860 29652
rect 27804 29598 27806 29650
rect 27806 29598 27858 29650
rect 27858 29598 27860 29650
rect 27804 29596 27860 29598
rect 27468 29484 27524 29540
rect 27916 29538 27972 29540
rect 27916 29486 27918 29538
rect 27918 29486 27970 29538
rect 27970 29486 27972 29538
rect 27916 29484 27972 29486
rect 27580 28812 27636 28868
rect 28588 30210 28644 30212
rect 28588 30158 28590 30210
rect 28590 30158 28642 30210
rect 28642 30158 28644 30210
rect 28588 30156 28644 30158
rect 28140 30098 28196 30100
rect 28140 30046 28142 30098
rect 28142 30046 28194 30098
rect 28194 30046 28196 30098
rect 28140 30044 28196 30046
rect 28588 29538 28644 29540
rect 28588 29486 28590 29538
rect 28590 29486 28642 29538
rect 28642 29486 28644 29538
rect 28588 29484 28644 29486
rect 28364 29426 28420 29428
rect 28364 29374 28366 29426
rect 28366 29374 28418 29426
rect 28418 29374 28420 29426
rect 28364 29372 28420 29374
rect 28700 29036 28756 29092
rect 29708 36482 29764 36484
rect 29708 36430 29710 36482
rect 29710 36430 29762 36482
rect 29762 36430 29764 36482
rect 29708 36428 29764 36430
rect 29820 34802 29876 34804
rect 29820 34750 29822 34802
rect 29822 34750 29874 34802
rect 29874 34750 29876 34802
rect 29820 34748 29876 34750
rect 30044 38162 30100 38164
rect 30044 38110 30046 38162
rect 30046 38110 30098 38162
rect 30098 38110 30100 38162
rect 30044 38108 30100 38110
rect 30044 37100 30100 37156
rect 30156 35868 30212 35924
rect 30044 34748 30100 34804
rect 30156 34690 30212 34692
rect 30156 34638 30158 34690
rect 30158 34638 30210 34690
rect 30210 34638 30212 34690
rect 30156 34636 30212 34638
rect 29932 34018 29988 34020
rect 29932 33966 29934 34018
rect 29934 33966 29986 34018
rect 29986 33966 29988 34018
rect 29932 33964 29988 33966
rect 29708 31554 29764 31556
rect 29708 31502 29710 31554
rect 29710 31502 29762 31554
rect 29762 31502 29764 31554
rect 29708 31500 29764 31502
rect 29708 31164 29764 31220
rect 29484 30994 29540 30996
rect 29484 30942 29486 30994
rect 29486 30942 29538 30994
rect 29538 30942 29540 30994
rect 29484 30940 29540 30942
rect 29036 29372 29092 29428
rect 28812 28812 28868 28868
rect 27468 28588 27524 28644
rect 29260 28700 29316 28756
rect 27580 28476 27636 28532
rect 27356 27970 27412 27972
rect 27356 27918 27358 27970
rect 27358 27918 27410 27970
rect 27410 27918 27412 27970
rect 27356 27916 27412 27918
rect 26684 27634 26740 27636
rect 26684 27582 26686 27634
rect 26686 27582 26738 27634
rect 26738 27582 26740 27634
rect 26684 27580 26740 27582
rect 28364 28588 28420 28644
rect 27020 26572 27076 26628
rect 28588 28642 28644 28644
rect 28588 28590 28590 28642
rect 28590 28590 28642 28642
rect 28642 28590 28644 28642
rect 28588 28588 28644 28590
rect 29148 28642 29204 28644
rect 29148 28590 29150 28642
rect 29150 28590 29202 28642
rect 29202 28590 29204 28642
rect 29148 28588 29204 28590
rect 25340 26348 25396 26404
rect 25228 26236 25284 26292
rect 25228 25900 25284 25956
rect 25228 25564 25284 25620
rect 27804 26348 27860 26404
rect 27132 25618 27188 25620
rect 27132 25566 27134 25618
rect 27134 25566 27186 25618
rect 27186 25566 27188 25618
rect 27132 25564 27188 25566
rect 27916 25506 27972 25508
rect 27916 25454 27918 25506
rect 27918 25454 27970 25506
rect 27970 25454 27972 25506
rect 27916 25452 27972 25454
rect 25004 24780 25060 24836
rect 24780 23938 24836 23940
rect 24780 23886 24782 23938
rect 24782 23886 24834 23938
rect 24834 23886 24836 23938
rect 24780 23884 24836 23886
rect 24556 23772 24612 23828
rect 25228 23772 25284 23828
rect 25788 24556 25844 24612
rect 26236 24610 26292 24612
rect 26236 24558 26238 24610
rect 26238 24558 26290 24610
rect 26290 24558 26292 24610
rect 26236 24556 26292 24558
rect 27916 24220 27972 24276
rect 25788 24050 25844 24052
rect 25788 23998 25790 24050
rect 25790 23998 25842 24050
rect 25842 23998 25844 24050
rect 25788 23996 25844 23998
rect 25452 23884 25508 23940
rect 22204 23266 22260 23268
rect 22204 23214 22206 23266
rect 22206 23214 22258 23266
rect 22258 23214 22260 23266
rect 22204 23212 22260 23214
rect 22988 23212 23044 23268
rect 28252 27916 28308 27972
rect 28140 27858 28196 27860
rect 28140 27806 28142 27858
rect 28142 27806 28194 27858
rect 28194 27806 28196 27858
rect 28140 27804 28196 27806
rect 29484 29036 29540 29092
rect 29596 28588 29652 28644
rect 29708 29372 29764 29428
rect 30380 39340 30436 39396
rect 30940 41804 30996 41860
rect 31388 41186 31444 41188
rect 31388 41134 31390 41186
rect 31390 41134 31442 41186
rect 31442 41134 31444 41186
rect 31388 41132 31444 41134
rect 31164 41074 31220 41076
rect 31164 41022 31166 41074
rect 31166 41022 31218 41074
rect 31218 41022 31220 41074
rect 31164 41020 31220 41022
rect 30828 40012 30884 40068
rect 30492 38556 30548 38612
rect 32060 47570 32116 47572
rect 32060 47518 32062 47570
rect 32062 47518 32114 47570
rect 32114 47518 32116 47570
rect 32060 47516 32116 47518
rect 31948 46732 32004 46788
rect 31836 45890 31892 45892
rect 31836 45838 31838 45890
rect 31838 45838 31890 45890
rect 31890 45838 31892 45890
rect 31836 45836 31892 45838
rect 31724 43650 31780 43652
rect 31724 43598 31726 43650
rect 31726 43598 31778 43650
rect 31778 43598 31780 43650
rect 31724 43596 31780 43598
rect 31724 39004 31780 39060
rect 31164 38668 31220 38724
rect 30604 37938 30660 37940
rect 30604 37886 30606 37938
rect 30606 37886 30658 37938
rect 30658 37886 30660 37938
rect 30604 37884 30660 37886
rect 30492 37042 30548 37044
rect 30492 36990 30494 37042
rect 30494 36990 30546 37042
rect 30546 36990 30548 37042
rect 30492 36988 30548 36990
rect 30380 34860 30436 34916
rect 30604 35308 30660 35364
rect 30380 34636 30436 34692
rect 30268 33516 30324 33572
rect 30492 33852 30548 33908
rect 30380 29596 30436 29652
rect 31052 38556 31108 38612
rect 31388 38444 31444 38500
rect 31164 38332 31220 38388
rect 30828 35196 30884 35252
rect 31052 34860 31108 34916
rect 30940 34690 30996 34692
rect 30940 34638 30942 34690
rect 30942 34638 30994 34690
rect 30994 34638 30996 34690
rect 30940 34636 30996 34638
rect 30940 33122 30996 33124
rect 30940 33070 30942 33122
rect 30942 33070 30994 33122
rect 30994 33070 30996 33122
rect 30940 33068 30996 33070
rect 30940 31554 30996 31556
rect 30940 31502 30942 31554
rect 30942 31502 30994 31554
rect 30994 31502 30996 31554
rect 30940 31500 30996 31502
rect 30940 30210 30996 30212
rect 30940 30158 30942 30210
rect 30942 30158 30994 30210
rect 30994 30158 30996 30210
rect 30940 30156 30996 30158
rect 30716 29932 30772 29988
rect 30492 28924 30548 28980
rect 31052 28252 31108 28308
rect 31276 38108 31332 38164
rect 32060 46002 32116 46004
rect 32060 45950 32062 46002
rect 32062 45950 32114 46002
rect 32114 45950 32116 46002
rect 32060 45948 32116 45950
rect 32172 45276 32228 45332
rect 32508 46956 32564 47012
rect 36092 54402 36148 54404
rect 36092 54350 36094 54402
rect 36094 54350 36146 54402
rect 36146 54350 36148 54402
rect 36092 54348 36148 54350
rect 38892 55804 38948 55860
rect 43260 56252 43316 56308
rect 44604 56306 44660 56308
rect 44604 56254 44606 56306
rect 44606 56254 44658 56306
rect 44658 56254 44660 56306
rect 44604 56252 44660 56254
rect 40460 55804 40516 55860
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 36876 54572 36932 54628
rect 36764 53676 36820 53732
rect 36540 53058 36596 53060
rect 36540 53006 36542 53058
rect 36542 53006 36594 53058
rect 36594 53006 36596 53058
rect 36540 53004 36596 53006
rect 35980 52780 36036 52836
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34860 52108 34916 52164
rect 36204 52274 36260 52276
rect 36204 52222 36206 52274
rect 36206 52222 36258 52274
rect 36258 52222 36260 52274
rect 36204 52220 36260 52222
rect 36316 52444 36372 52500
rect 35980 52108 36036 52164
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 33180 50034 33236 50036
rect 33180 49982 33182 50034
rect 33182 49982 33234 50034
rect 33234 49982 33236 50034
rect 33180 49980 33236 49982
rect 32844 49196 32900 49252
rect 34188 49196 34244 49252
rect 32620 46396 32676 46452
rect 33068 49084 33124 49140
rect 34300 49026 34356 49028
rect 34300 48974 34302 49026
rect 34302 48974 34354 49026
rect 34354 48974 34356 49026
rect 34300 48972 34356 48974
rect 32956 48802 33012 48804
rect 32956 48750 32958 48802
rect 32958 48750 33010 48802
rect 33010 48750 33012 48802
rect 32956 48748 33012 48750
rect 33292 48802 33348 48804
rect 33292 48750 33294 48802
rect 33294 48750 33346 48802
rect 33346 48750 33348 48802
rect 33292 48748 33348 48750
rect 33068 48524 33124 48580
rect 33068 47404 33124 47460
rect 32956 46060 33012 46116
rect 33516 47964 33572 48020
rect 33852 47628 33908 47684
rect 33740 47458 33796 47460
rect 33740 47406 33742 47458
rect 33742 47406 33794 47458
rect 33794 47406 33796 47458
rect 33740 47404 33796 47406
rect 33628 46956 33684 47012
rect 34636 48802 34692 48804
rect 34636 48750 34638 48802
rect 34638 48750 34690 48802
rect 34690 48750 34692 48802
rect 34636 48748 34692 48750
rect 34860 47628 34916 47684
rect 34188 47180 34244 47236
rect 33740 47068 33796 47124
rect 33180 45778 33236 45780
rect 33180 45726 33182 45778
rect 33182 45726 33234 45778
rect 33234 45726 33236 45778
rect 33180 45724 33236 45726
rect 34076 46898 34132 46900
rect 34076 46846 34078 46898
rect 34078 46846 34130 46898
rect 34130 46846 34132 46898
rect 34076 46844 34132 46846
rect 33292 46396 33348 46452
rect 32732 45612 32788 45668
rect 32508 45106 32564 45108
rect 32508 45054 32510 45106
rect 32510 45054 32562 45106
rect 32562 45054 32564 45106
rect 32508 45052 32564 45054
rect 32396 44492 32452 44548
rect 32060 44044 32116 44100
rect 32508 43426 32564 43428
rect 32508 43374 32510 43426
rect 32510 43374 32562 43426
rect 32562 43374 32564 43426
rect 32508 43372 32564 43374
rect 32060 41916 32116 41972
rect 33404 45106 33460 45108
rect 33404 45054 33406 45106
rect 33406 45054 33458 45106
rect 33458 45054 33460 45106
rect 33404 45052 33460 45054
rect 33852 44492 33908 44548
rect 33516 44434 33572 44436
rect 33516 44382 33518 44434
rect 33518 44382 33570 44434
rect 33570 44382 33572 44434
rect 33516 44380 33572 44382
rect 33068 42812 33124 42868
rect 34524 46562 34580 46564
rect 34524 46510 34526 46562
rect 34526 46510 34578 46562
rect 34578 46510 34580 46562
rect 34524 46508 34580 46510
rect 34748 45778 34804 45780
rect 34748 45726 34750 45778
rect 34750 45726 34802 45778
rect 34802 45726 34804 45778
rect 34748 45724 34804 45726
rect 34300 45666 34356 45668
rect 34300 45614 34302 45666
rect 34302 45614 34354 45666
rect 34354 45614 34356 45666
rect 34300 45612 34356 45614
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35084 49026 35140 49028
rect 35084 48974 35086 49026
rect 35086 48974 35138 49026
rect 35138 48974 35140 49026
rect 35084 48972 35140 48974
rect 35420 49026 35476 49028
rect 35420 48974 35422 49026
rect 35422 48974 35474 49026
rect 35474 48974 35476 49026
rect 35420 48972 35476 48974
rect 35980 48972 36036 49028
rect 35644 48412 35700 48468
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35644 47628 35700 47684
rect 35196 47068 35252 47124
rect 35084 46732 35140 46788
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35644 45612 35700 45668
rect 35644 45276 35700 45332
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 33964 43708 34020 43764
rect 33404 43650 33460 43652
rect 33404 43598 33406 43650
rect 33406 43598 33458 43650
rect 33458 43598 33460 43650
rect 33404 43596 33460 43598
rect 33292 43484 33348 43540
rect 33180 43372 33236 43428
rect 33516 43260 33572 43316
rect 33852 42924 33908 42980
rect 34748 44322 34804 44324
rect 34748 44270 34750 44322
rect 34750 44270 34802 44322
rect 34802 44270 34804 44322
rect 34748 44268 34804 44270
rect 35420 44268 35476 44324
rect 34972 43596 35028 43652
rect 34748 42866 34804 42868
rect 34748 42814 34750 42866
rect 34750 42814 34802 42866
rect 34802 42814 34804 42866
rect 34748 42812 34804 42814
rect 34524 42252 34580 42308
rect 33964 41970 34020 41972
rect 33964 41918 33966 41970
rect 33966 41918 34018 41970
rect 34018 41918 34020 41970
rect 33964 41916 34020 41918
rect 33852 41692 33908 41748
rect 32956 40962 33012 40964
rect 32956 40910 32958 40962
rect 32958 40910 33010 40962
rect 33010 40910 33012 40962
rect 32956 40908 33012 40910
rect 32172 40796 32228 40852
rect 34524 41916 34580 41972
rect 32284 40348 32340 40404
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35308 42812 35364 42868
rect 34524 40796 34580 40852
rect 34636 41132 34692 41188
rect 35420 42252 35476 42308
rect 37100 52892 37156 52948
rect 36988 52274 37044 52276
rect 36988 52222 36990 52274
rect 36990 52222 37042 52274
rect 37042 52222 37044 52274
rect 36988 52220 37044 52222
rect 37660 53900 37716 53956
rect 38108 54684 38164 54740
rect 38220 54514 38276 54516
rect 38220 54462 38222 54514
rect 38222 54462 38274 54514
rect 38274 54462 38276 54514
rect 38220 54460 38276 54462
rect 38108 53900 38164 53956
rect 38556 54514 38612 54516
rect 38556 54462 38558 54514
rect 38558 54462 38610 54514
rect 38610 54462 38612 54514
rect 38556 54460 38612 54462
rect 38892 54460 38948 54516
rect 39900 55074 39956 55076
rect 39900 55022 39902 55074
rect 39902 55022 39954 55074
rect 39954 55022 39956 55074
rect 39900 55020 39956 55022
rect 40236 55020 40292 55076
rect 41916 55020 41972 55076
rect 39564 54626 39620 54628
rect 39564 54574 39566 54626
rect 39566 54574 39618 54626
rect 39618 54574 39620 54626
rect 39564 54572 39620 54574
rect 40908 54626 40964 54628
rect 40908 54574 40910 54626
rect 40910 54574 40962 54626
rect 40962 54574 40964 54626
rect 40908 54572 40964 54574
rect 39004 54348 39060 54404
rect 38220 53788 38276 53844
rect 38780 54012 38836 54068
rect 37324 52444 37380 52500
rect 37212 52108 37268 52164
rect 37324 51660 37380 51716
rect 38668 52332 38724 52388
rect 38220 52162 38276 52164
rect 38220 52110 38222 52162
rect 38222 52110 38274 52162
rect 38274 52110 38276 52162
rect 38220 52108 38276 52110
rect 38108 51660 38164 51716
rect 37996 51548 38052 51604
rect 40348 54402 40404 54404
rect 40348 54350 40350 54402
rect 40350 54350 40402 54402
rect 40402 54350 40404 54402
rect 40348 54348 40404 54350
rect 38892 53842 38948 53844
rect 38892 53790 38894 53842
rect 38894 53790 38946 53842
rect 38946 53790 38948 53842
rect 38892 53788 38948 53790
rect 41356 54514 41412 54516
rect 41356 54462 41358 54514
rect 41358 54462 41410 54514
rect 41410 54462 41412 54514
rect 41356 54460 41412 54462
rect 41132 54348 41188 54404
rect 40908 53954 40964 53956
rect 40908 53902 40910 53954
rect 40910 53902 40962 53954
rect 40962 53902 40964 53954
rect 40908 53900 40964 53902
rect 41580 54460 41636 54516
rect 41244 53730 41300 53732
rect 41244 53678 41246 53730
rect 41246 53678 41298 53730
rect 41298 53678 41300 53730
rect 41244 53676 41300 53678
rect 40348 52834 40404 52836
rect 40348 52782 40350 52834
rect 40350 52782 40402 52834
rect 40402 52782 40404 52834
rect 40348 52780 40404 52782
rect 39116 52050 39172 52052
rect 39116 51998 39118 52050
rect 39118 51998 39170 52050
rect 39170 51998 39172 52050
rect 39116 51996 39172 51998
rect 38892 51602 38948 51604
rect 38892 51550 38894 51602
rect 38894 51550 38946 51602
rect 38946 51550 38948 51602
rect 38892 51548 38948 51550
rect 40124 51602 40180 51604
rect 40124 51550 40126 51602
rect 40126 51550 40178 51602
rect 40178 51550 40180 51602
rect 40124 51548 40180 51550
rect 39676 51490 39732 51492
rect 39676 51438 39678 51490
rect 39678 51438 39730 51490
rect 39730 51438 39732 51490
rect 39676 51436 39732 51438
rect 38556 51266 38612 51268
rect 38556 51214 38558 51266
rect 38558 51214 38610 51266
rect 38610 51214 38612 51266
rect 38556 51212 38612 51214
rect 36428 50594 36484 50596
rect 36428 50542 36430 50594
rect 36430 50542 36482 50594
rect 36482 50542 36484 50594
rect 36428 50540 36484 50542
rect 37324 50594 37380 50596
rect 37324 50542 37326 50594
rect 37326 50542 37378 50594
rect 37378 50542 37380 50594
rect 37324 50540 37380 50542
rect 38444 49868 38500 49924
rect 36316 48412 36372 48468
rect 38220 48130 38276 48132
rect 38220 48078 38222 48130
rect 38222 48078 38274 48130
rect 38274 48078 38276 48130
rect 38220 48076 38276 48078
rect 38108 47458 38164 47460
rect 38108 47406 38110 47458
rect 38110 47406 38162 47458
rect 38162 47406 38164 47458
rect 38108 47404 38164 47406
rect 39228 51154 39284 51156
rect 39228 51102 39230 51154
rect 39230 51102 39282 51154
rect 39282 51102 39284 51154
rect 39228 51100 39284 51102
rect 39452 51378 39508 51380
rect 39452 51326 39454 51378
rect 39454 51326 39506 51378
rect 39506 51326 39508 51378
rect 39452 51324 39508 51326
rect 41132 52780 41188 52836
rect 41356 53170 41412 53172
rect 41356 53118 41358 53170
rect 41358 53118 41410 53170
rect 41410 53118 41412 53170
rect 41356 53116 41412 53118
rect 41692 53788 41748 53844
rect 42028 53842 42084 53844
rect 42028 53790 42030 53842
rect 42030 53790 42082 53842
rect 42082 53790 42084 53842
rect 42028 53788 42084 53790
rect 47740 56252 47796 56308
rect 48972 56306 49028 56308
rect 48972 56254 48974 56306
rect 48974 56254 49026 56306
rect 49026 56254 49028 56306
rect 48972 56252 49028 56254
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 49980 56252 50036 56308
rect 52220 56306 52276 56308
rect 52220 56254 52222 56306
rect 52222 56254 52274 56306
rect 52274 56254 52276 56306
rect 52220 56252 52276 56254
rect 45500 55356 45556 55412
rect 46732 55410 46788 55412
rect 46732 55358 46734 55410
rect 46734 55358 46786 55410
rect 46786 55358 46788 55410
rect 46732 55356 46788 55358
rect 43484 54012 43540 54068
rect 42924 53676 42980 53732
rect 41244 52444 41300 52500
rect 40908 51436 40964 51492
rect 40348 51212 40404 51268
rect 38892 48300 38948 48356
rect 38556 47458 38612 47460
rect 38556 47406 38558 47458
rect 38558 47406 38610 47458
rect 38610 47406 38612 47458
rect 38556 47404 38612 47406
rect 36652 46786 36708 46788
rect 36652 46734 36654 46786
rect 36654 46734 36706 46786
rect 36706 46734 36708 46786
rect 36652 46732 36708 46734
rect 38780 46956 38836 47012
rect 38444 46508 38500 46564
rect 38668 45836 38724 45892
rect 38668 45666 38724 45668
rect 38668 45614 38670 45666
rect 38670 45614 38722 45666
rect 38722 45614 38724 45666
rect 38668 45612 38724 45614
rect 36204 44492 36260 44548
rect 37100 44268 37156 44324
rect 37100 43708 37156 43764
rect 35980 42700 36036 42756
rect 35532 41916 35588 41972
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 41020 35252 41076
rect 36316 41858 36372 41860
rect 36316 41806 36318 41858
rect 36318 41806 36370 41858
rect 36370 41806 36372 41858
rect 36316 41804 36372 41806
rect 35420 41186 35476 41188
rect 35420 41134 35422 41186
rect 35422 41134 35474 41186
rect 35474 41134 35476 41186
rect 35420 41132 35476 41134
rect 35308 40572 35364 40628
rect 34748 40348 34804 40404
rect 35532 40402 35588 40404
rect 35532 40350 35534 40402
rect 35534 40350 35586 40402
rect 35586 40350 35588 40402
rect 35532 40348 35588 40350
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 31948 38780 32004 38836
rect 32060 37938 32116 37940
rect 32060 37886 32062 37938
rect 32062 37886 32114 37938
rect 32114 37886 32116 37938
rect 32060 37884 32116 37886
rect 31724 37772 31780 37828
rect 32172 37772 32228 37828
rect 32508 38556 32564 38612
rect 32956 38556 33012 38612
rect 32396 38444 32452 38500
rect 31500 37324 31556 37380
rect 33628 38780 33684 38836
rect 33852 38722 33908 38724
rect 33852 38670 33854 38722
rect 33854 38670 33906 38722
rect 33906 38670 33908 38722
rect 33852 38668 33908 38670
rect 33516 38556 33572 38612
rect 33404 37884 33460 37940
rect 33292 37772 33348 37828
rect 32060 37212 32116 37268
rect 31948 37154 32004 37156
rect 31948 37102 31950 37154
rect 31950 37102 32002 37154
rect 32002 37102 32004 37154
rect 31948 37100 32004 37102
rect 31388 35308 31444 35364
rect 31724 35644 31780 35700
rect 31724 34748 31780 34804
rect 31388 33068 31444 33124
rect 31500 30044 31556 30100
rect 32396 37212 32452 37268
rect 32956 37436 33012 37492
rect 32172 34860 32228 34916
rect 32508 33852 32564 33908
rect 32396 33740 32452 33796
rect 32396 33404 32452 33460
rect 33180 35196 33236 35252
rect 33068 34860 33124 34916
rect 33068 33740 33124 33796
rect 33516 35980 33572 36036
rect 33516 35308 33572 35364
rect 35644 39004 35700 39060
rect 35756 38892 35812 38948
rect 34188 38108 34244 38164
rect 33852 37826 33908 37828
rect 33852 37774 33854 37826
rect 33854 37774 33906 37826
rect 33906 37774 33908 37826
rect 33852 37772 33908 37774
rect 34300 37266 34356 37268
rect 34300 37214 34302 37266
rect 34302 37214 34354 37266
rect 34354 37214 34356 37266
rect 34300 37212 34356 37214
rect 34076 35644 34132 35700
rect 34188 35308 34244 35364
rect 34636 36594 34692 36596
rect 34636 36542 34638 36594
rect 34638 36542 34690 36594
rect 34690 36542 34692 36594
rect 34636 36540 34692 36542
rect 34748 35922 34804 35924
rect 34748 35870 34750 35922
rect 34750 35870 34802 35922
rect 34802 35870 34804 35922
rect 34748 35868 34804 35870
rect 34860 35756 34916 35812
rect 34748 35308 34804 35364
rect 34636 34690 34692 34692
rect 34636 34638 34638 34690
rect 34638 34638 34690 34690
rect 34690 34638 34692 34690
rect 34636 34636 34692 34638
rect 33404 33404 33460 33460
rect 33516 33516 33572 33572
rect 32060 31836 32116 31892
rect 32396 31836 32452 31892
rect 33068 31836 33124 31892
rect 33628 32674 33684 32676
rect 33628 32622 33630 32674
rect 33630 32622 33682 32674
rect 33682 32622 33684 32674
rect 33628 32620 33684 32622
rect 33964 32620 34020 32676
rect 33180 31218 33236 31220
rect 33180 31166 33182 31218
rect 33182 31166 33234 31218
rect 33234 31166 33236 31218
rect 33180 31164 33236 31166
rect 33964 30940 34020 30996
rect 35532 38668 35588 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 36204 40796 36260 40852
rect 36316 40626 36372 40628
rect 36316 40574 36318 40626
rect 36318 40574 36370 40626
rect 36370 40574 36372 40626
rect 36316 40572 36372 40574
rect 36764 40460 36820 40516
rect 36876 42700 36932 42756
rect 36876 41020 36932 41076
rect 37212 43596 37268 43652
rect 37436 44156 37492 44212
rect 38780 43650 38836 43652
rect 38780 43598 38782 43650
rect 38782 43598 38834 43650
rect 38834 43598 38836 43650
rect 38780 43596 38836 43598
rect 39116 46508 39172 46564
rect 39676 48130 39732 48132
rect 39676 48078 39678 48130
rect 39678 48078 39730 48130
rect 39730 48078 39732 48130
rect 39676 48076 39732 48078
rect 39452 46956 39508 47012
rect 39228 46620 39284 46676
rect 39564 46732 39620 46788
rect 40908 50594 40964 50596
rect 40908 50542 40910 50594
rect 40910 50542 40962 50594
rect 40962 50542 40964 50594
rect 40908 50540 40964 50542
rect 41468 51100 41524 51156
rect 42140 52050 42196 52052
rect 42140 51998 42142 52050
rect 42142 51998 42194 52050
rect 42194 51998 42196 52050
rect 42140 51996 42196 51998
rect 41132 50428 41188 50484
rect 40908 46786 40964 46788
rect 40908 46734 40910 46786
rect 40910 46734 40962 46786
rect 40962 46734 40964 46786
rect 40908 46732 40964 46734
rect 39228 45612 39284 45668
rect 40236 46620 40292 46676
rect 40012 44322 40068 44324
rect 40012 44270 40014 44322
rect 40014 44270 40066 44322
rect 40066 44270 40068 44322
rect 40012 44268 40068 44270
rect 39676 43708 39732 43764
rect 37324 43538 37380 43540
rect 37324 43486 37326 43538
rect 37326 43486 37378 43538
rect 37378 43486 37380 43538
rect 37324 43484 37380 43486
rect 39452 43650 39508 43652
rect 39452 43598 39454 43650
rect 39454 43598 39506 43650
rect 39506 43598 39508 43650
rect 39452 43596 39508 43598
rect 39228 43484 39284 43540
rect 38668 43314 38724 43316
rect 38668 43262 38670 43314
rect 38670 43262 38722 43314
rect 38722 43262 38724 43314
rect 38668 43260 38724 43262
rect 40124 42754 40180 42756
rect 40124 42702 40126 42754
rect 40126 42702 40178 42754
rect 40178 42702 40180 42754
rect 40124 42700 40180 42702
rect 42812 53116 42868 53172
rect 42588 52780 42644 52836
rect 42252 51602 42308 51604
rect 42252 51550 42254 51602
rect 42254 51550 42306 51602
rect 42306 51550 42308 51602
rect 42252 51548 42308 51550
rect 44604 53788 44660 53844
rect 42476 50652 42532 50708
rect 44156 50706 44212 50708
rect 44156 50654 44158 50706
rect 44158 50654 44210 50706
rect 44210 50654 44212 50706
rect 44156 50652 44212 50654
rect 41356 50594 41412 50596
rect 41356 50542 41358 50594
rect 41358 50542 41410 50594
rect 41410 50542 41412 50594
rect 41356 50540 41412 50542
rect 42028 50482 42084 50484
rect 42028 50430 42030 50482
rect 42030 50430 42082 50482
rect 42082 50430 42084 50482
rect 42028 50428 42084 50430
rect 42812 48076 42868 48132
rect 41356 47292 41412 47348
rect 42140 47346 42196 47348
rect 42140 47294 42142 47346
rect 42142 47294 42194 47346
rect 42194 47294 42196 47346
rect 42140 47292 42196 47294
rect 41468 46674 41524 46676
rect 41468 46622 41470 46674
rect 41470 46622 41522 46674
rect 41522 46622 41524 46674
rect 41468 46620 41524 46622
rect 41020 45276 41076 45332
rect 41020 44940 41076 44996
rect 40572 43596 40628 43652
rect 40908 44268 40964 44324
rect 40684 42754 40740 42756
rect 40684 42702 40686 42754
rect 40686 42702 40738 42754
rect 40738 42702 40740 42754
rect 40684 42700 40740 42702
rect 37772 41916 37828 41972
rect 40124 41858 40180 41860
rect 40124 41806 40126 41858
rect 40126 41806 40178 41858
rect 40178 41806 40180 41858
rect 40124 41804 40180 41806
rect 40012 41746 40068 41748
rect 40012 41694 40014 41746
rect 40014 41694 40066 41746
rect 40066 41694 40068 41746
rect 40012 41692 40068 41694
rect 44492 44994 44548 44996
rect 44492 44942 44494 44994
rect 44494 44942 44546 44994
rect 44546 44942 44548 44994
rect 44492 44940 44548 44942
rect 41580 44268 41636 44324
rect 41020 44156 41076 44212
rect 41132 43762 41188 43764
rect 41132 43710 41134 43762
rect 41134 43710 41186 43762
rect 41186 43710 41188 43762
rect 41132 43708 41188 43710
rect 41580 43650 41636 43652
rect 41580 43598 41582 43650
rect 41582 43598 41634 43650
rect 41634 43598 41636 43650
rect 41580 43596 41636 43598
rect 44940 52834 44996 52836
rect 44940 52782 44942 52834
rect 44942 52782 44994 52834
rect 44994 52782 44996 52834
rect 44940 52780 44996 52782
rect 45388 48972 45444 49028
rect 54460 56252 54516 56308
rect 56028 56306 56084 56308
rect 56028 56254 56030 56306
rect 56030 56254 56082 56306
rect 56082 56254 56084 56306
rect 56028 56252 56084 56254
rect 52332 55356 52388 55412
rect 53676 55410 53732 55412
rect 53676 55358 53678 55410
rect 53678 55358 53730 55410
rect 53730 55358 53732 55410
rect 53676 55356 53732 55358
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 47740 47516 47796 47572
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50316 45948 50372 46004
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 44604 42924 44660 42980
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 41356 41916 41412 41972
rect 43820 41858 43876 41860
rect 43820 41806 43822 41858
rect 43822 41806 43874 41858
rect 43874 41806 43876 41858
rect 43820 41804 43876 41806
rect 36428 39004 36484 39060
rect 36092 37212 36148 37268
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36316 36876 36372 36932
rect 36092 36540 36148 36596
rect 35532 35980 35588 36036
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35084 34914 35140 34916
rect 35084 34862 35086 34914
rect 35086 34862 35138 34914
rect 35138 34862 35140 34914
rect 35084 34860 35140 34862
rect 38444 40460 38500 40516
rect 38220 38946 38276 38948
rect 38220 38894 38222 38946
rect 38222 38894 38274 38946
rect 38274 38894 38276 38946
rect 38220 38892 38276 38894
rect 36988 38668 37044 38724
rect 37436 38668 37492 38724
rect 37772 38668 37828 38724
rect 37212 38220 37268 38276
rect 36764 36876 36820 36932
rect 36652 36540 36708 36596
rect 36316 36482 36372 36484
rect 36316 36430 36318 36482
rect 36318 36430 36370 36482
rect 36370 36430 36372 36482
rect 36316 36428 36372 36430
rect 37324 35756 37380 35812
rect 36428 35308 36484 35364
rect 34972 34412 35028 34468
rect 36316 34524 36372 34580
rect 34412 34130 34468 34132
rect 34412 34078 34414 34130
rect 34414 34078 34466 34130
rect 34466 34078 34468 34130
rect 34412 34076 34468 34078
rect 34300 33516 34356 33572
rect 34076 31052 34132 31108
rect 34188 33404 34244 33460
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34748 33516 34804 33572
rect 34524 31724 34580 31780
rect 31948 30210 32004 30212
rect 31948 30158 31950 30210
rect 31950 30158 32002 30210
rect 32002 30158 32004 30210
rect 31948 30156 32004 30158
rect 35308 33122 35364 33124
rect 35308 33070 35310 33122
rect 35310 33070 35362 33122
rect 35362 33070 35364 33122
rect 35308 33068 35364 33070
rect 35868 33852 35924 33908
rect 37660 35980 37716 36036
rect 37772 35810 37828 35812
rect 37772 35758 37774 35810
rect 37774 35758 37826 35810
rect 37826 35758 37828 35810
rect 37772 35756 37828 35758
rect 37548 35308 37604 35364
rect 37548 34748 37604 34804
rect 37436 34524 37492 34580
rect 36652 34130 36708 34132
rect 36652 34078 36654 34130
rect 36654 34078 36706 34130
rect 36706 34078 36708 34130
rect 36652 34076 36708 34078
rect 34636 30156 34692 30212
rect 35756 32396 35812 32452
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 37100 33852 37156 33908
rect 37100 33346 37156 33348
rect 37100 33294 37102 33346
rect 37102 33294 37154 33346
rect 37154 33294 37156 33346
rect 37100 33292 37156 33294
rect 38220 37436 38276 37492
rect 54572 53788 54628 53844
rect 55356 44380 55412 44436
rect 52668 40908 52724 40964
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 39900 38668 39956 38724
rect 38108 35868 38164 35924
rect 37772 33292 37828 33348
rect 39564 37490 39620 37492
rect 39564 37438 39566 37490
rect 39566 37438 39618 37490
rect 39618 37438 39620 37490
rect 39564 37436 39620 37438
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 38892 36428 38948 36484
rect 38220 34300 38276 34356
rect 38668 35868 38724 35924
rect 37212 33122 37268 33124
rect 37212 33070 37214 33122
rect 37214 33070 37266 33122
rect 37266 33070 37268 33122
rect 37212 33068 37268 33070
rect 37548 32450 37604 32452
rect 37548 32398 37550 32450
rect 37550 32398 37602 32450
rect 37602 32398 37604 32450
rect 37548 32396 37604 32398
rect 36092 31666 36148 31668
rect 36092 31614 36094 31666
rect 36094 31614 36146 31666
rect 36146 31614 36148 31666
rect 36092 31612 36148 31614
rect 35756 31106 35812 31108
rect 35756 31054 35758 31106
rect 35758 31054 35810 31106
rect 35810 31054 35812 31106
rect 35756 31052 35812 31054
rect 35980 30940 36036 30996
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34860 30210 34916 30212
rect 34860 30158 34862 30210
rect 34862 30158 34914 30210
rect 34914 30158 34916 30210
rect 34860 30156 34916 30158
rect 35868 30210 35924 30212
rect 35868 30158 35870 30210
rect 35870 30158 35922 30210
rect 35922 30158 35924 30210
rect 35868 30156 35924 30158
rect 31836 29148 31892 29204
rect 31164 28140 31220 28196
rect 29932 28082 29988 28084
rect 29932 28030 29934 28082
rect 29934 28030 29986 28082
rect 29986 28030 29988 28082
rect 29932 28028 29988 28030
rect 30828 28082 30884 28084
rect 30828 28030 30830 28082
rect 30830 28030 30882 28082
rect 30882 28030 30884 28082
rect 30828 28028 30884 28030
rect 30268 27970 30324 27972
rect 30268 27918 30270 27970
rect 30270 27918 30322 27970
rect 30322 27918 30324 27970
rect 30268 27916 30324 27918
rect 29260 27468 29316 27524
rect 28252 26348 28308 26404
rect 29260 25452 29316 25508
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 36988 31778 37044 31780
rect 36988 31726 36990 31778
rect 36990 31726 37042 31778
rect 37042 31726 37044 31778
rect 36988 31724 37044 31726
rect 37884 31724 37940 31780
rect 36876 30994 36932 30996
rect 36876 30942 36878 30994
rect 36878 30942 36930 30994
rect 36930 30942 36932 30994
rect 36876 30940 36932 30942
rect 36204 30322 36260 30324
rect 36204 30270 36206 30322
rect 36206 30270 36258 30322
rect 36258 30270 36260 30322
rect 36204 30268 36260 30270
rect 37324 31612 37380 31668
rect 37212 31554 37268 31556
rect 37212 31502 37214 31554
rect 37214 31502 37266 31554
rect 37266 31502 37268 31554
rect 37212 31500 37268 31502
rect 36988 30156 37044 30212
rect 39340 35922 39396 35924
rect 39340 35870 39342 35922
rect 39342 35870 39394 35922
rect 39394 35870 39396 35922
rect 39340 35868 39396 35870
rect 39228 34354 39284 34356
rect 39228 34302 39230 34354
rect 39230 34302 39282 34354
rect 39282 34302 39284 34354
rect 39228 34300 39284 34302
rect 39340 34188 39396 34244
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 39788 34188 39844 34244
rect 39900 35308 39956 35364
rect 40012 33516 40068 33572
rect 38332 33068 38388 33124
rect 38220 30268 38276 30324
rect 35644 28028 35700 28084
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34860 25564 34916 25620
rect 29372 25116 29428 25172
rect 39564 32620 39620 32676
rect 41916 34524 41972 34580
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 41468 33516 41524 33572
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 39116 31778 39172 31780
rect 39116 31726 39118 31778
rect 39118 31726 39170 31778
rect 39170 31726 39172 31778
rect 39116 31724 39172 31726
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 39004 24556 39060 24612
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 28028 22876 28084 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 6748 9660 6804 9716
rect 5628 9436 5684 9492
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 5068 6748 5124 6804
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 2492 3836 2548 3892
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 1708 3276 1764 3332
rect 2716 3276 2772 3332
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 1708 2044 1764 2100
<< metal3 >>
rect 0 57652 800 57680
rect 0 57596 2156 57652
rect 2212 57596 2222 57652
rect 0 57568 800 57596
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 43250 56252 43260 56308
rect 43316 56252 44604 56308
rect 44660 56252 44670 56308
rect 47730 56252 47740 56308
rect 47796 56252 48972 56308
rect 49028 56252 49038 56308
rect 49970 56252 49980 56308
rect 50036 56252 52220 56308
rect 52276 56252 52286 56308
rect 54450 56252 54460 56308
rect 54516 56252 56028 56308
rect 56084 56252 56094 56308
rect 2146 56028 2156 56084
rect 2212 56028 2604 56084
rect 2660 56028 2670 56084
rect 27906 55916 27916 55972
rect 27972 55916 28588 55972
rect 28644 55916 28654 55972
rect 0 55860 800 55888
rect 0 55804 1708 55860
rect 1764 55804 3164 55860
rect 3220 55804 3230 55860
rect 28354 55804 28364 55860
rect 28420 55804 38892 55860
rect 38948 55804 40460 55860
rect 40516 55804 40526 55860
rect 0 55776 800 55804
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 18498 55356 18508 55412
rect 18564 55356 20524 55412
rect 20580 55356 23324 55412
rect 23380 55356 23390 55412
rect 45490 55356 45500 55412
rect 45556 55356 46732 55412
rect 46788 55356 46798 55412
rect 52322 55356 52332 55412
rect 52388 55356 53676 55412
rect 53732 55356 53742 55412
rect 13570 55244 13580 55300
rect 13636 55244 16828 55300
rect 16884 55244 17724 55300
rect 17780 55244 18732 55300
rect 18788 55244 21420 55300
rect 21476 55244 21486 55300
rect 29250 55244 29260 55300
rect 29316 55244 33180 55300
rect 33236 55244 33246 55300
rect 5842 55132 5852 55188
rect 5908 55132 11788 55188
rect 11844 55132 11854 55188
rect 22642 55020 22652 55076
rect 22708 55020 27580 55076
rect 27636 55020 32508 55076
rect 32564 55020 32574 55076
rect 39890 55020 39900 55076
rect 39956 55020 40236 55076
rect 40292 55020 41916 55076
rect 41972 55020 41982 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 31892 54684 36092 54740
rect 36148 54684 38108 54740
rect 38164 54684 38174 54740
rect 1586 54572 1596 54628
rect 1652 54572 2044 54628
rect 2100 54572 2110 54628
rect 12338 54572 12348 54628
rect 12404 54572 29148 54628
rect 29204 54572 29214 54628
rect 31826 54572 31836 54628
rect 31892 54572 31948 54684
rect 32498 54572 32508 54628
rect 32564 54572 33404 54628
rect 33460 54572 33470 54628
rect 33618 54572 33628 54628
rect 33684 54572 36876 54628
rect 36932 54572 36942 54628
rect 39554 54572 39564 54628
rect 39620 54572 40908 54628
rect 40964 54572 40974 54628
rect 15698 54460 15708 54516
rect 15764 54460 16828 54516
rect 16884 54460 16894 54516
rect 17826 54460 17836 54516
rect 17892 54460 18396 54516
rect 18452 54460 18462 54516
rect 22866 54460 22876 54516
rect 22932 54460 23436 54516
rect 23492 54460 28812 54516
rect 28868 54460 30044 54516
rect 30100 54460 30110 54516
rect 33842 54460 33852 54516
rect 33908 54460 38220 54516
rect 38276 54460 38556 54516
rect 38612 54460 38622 54516
rect 38882 54460 38892 54516
rect 38948 54460 41356 54516
rect 41412 54460 41580 54516
rect 41636 54460 41646 54516
rect 16828 54404 16884 54460
rect 16828 54348 18284 54404
rect 18340 54348 18350 54404
rect 24770 54348 24780 54404
rect 24836 54348 26012 54404
rect 26068 54348 26078 54404
rect 33954 54348 33964 54404
rect 34020 54348 36092 54404
rect 36148 54348 36158 54404
rect 38994 54348 39004 54404
rect 39060 54348 40348 54404
rect 40404 54348 41132 54404
rect 41188 54348 41198 54404
rect 0 54068 800 54096
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 0 54012 1708 54068
rect 1764 54012 2492 54068
rect 2548 54012 2558 54068
rect 38770 54012 38780 54068
rect 38836 54012 43484 54068
rect 43540 54012 43550 54068
rect 0 53984 800 54012
rect 29250 53900 29260 53956
rect 29316 53900 37660 53956
rect 37716 53900 37726 53956
rect 38098 53900 38108 53956
rect 38164 53900 40908 53956
rect 40964 53900 40974 53956
rect 2930 53788 2940 53844
rect 2996 53788 5628 53844
rect 5684 53788 5694 53844
rect 15922 53788 15932 53844
rect 15988 53788 16604 53844
rect 16660 53788 18844 53844
rect 18900 53788 18910 53844
rect 21532 53788 21980 53844
rect 22036 53788 22652 53844
rect 22708 53788 22718 53844
rect 22866 53788 22876 53844
rect 22932 53788 23660 53844
rect 23716 53788 23726 53844
rect 25106 53788 25116 53844
rect 25172 53788 26348 53844
rect 26404 53788 26414 53844
rect 26562 53788 26572 53844
rect 26628 53788 28140 53844
rect 28196 53788 28206 53844
rect 30370 53788 30380 53844
rect 30436 53788 33292 53844
rect 33348 53788 33628 53844
rect 33684 53788 33694 53844
rect 38210 53788 38220 53844
rect 38276 53788 38892 53844
rect 38948 53788 38958 53844
rect 41682 53788 41692 53844
rect 41748 53788 42028 53844
rect 42084 53788 42094 53844
rect 44594 53788 44604 53844
rect 44660 53788 54572 53844
rect 54628 53788 54638 53844
rect 21532 53732 21588 53788
rect 17602 53676 17612 53732
rect 17668 53676 18172 53732
rect 18228 53676 21588 53732
rect 21746 53676 21756 53732
rect 21812 53676 22428 53732
rect 22484 53676 22494 53732
rect 32050 53676 32060 53732
rect 32116 53676 36764 53732
rect 36820 53676 36830 53732
rect 41234 53676 41244 53732
rect 41300 53676 42924 53732
rect 42980 53676 42990 53732
rect 12786 53564 12796 53620
rect 12852 53564 13804 53620
rect 13860 53564 32620 53620
rect 32676 53564 33068 53620
rect 33124 53564 33852 53620
rect 33908 53564 34636 53620
rect 34692 53564 34702 53620
rect 10882 53452 10892 53508
rect 10948 53452 11564 53508
rect 11620 53452 17612 53508
rect 17668 53452 17678 53508
rect 22306 53452 22316 53508
rect 22372 53452 24444 53508
rect 24500 53452 24510 53508
rect 24882 53452 24892 53508
rect 24948 53452 25564 53508
rect 25620 53452 29148 53508
rect 29204 53452 30156 53508
rect 30212 53452 30222 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 12898 53116 12908 53172
rect 12964 53116 15932 53172
rect 15988 53116 16380 53172
rect 16436 53116 27076 53172
rect 7970 53004 7980 53060
rect 8036 53004 10668 53060
rect 10724 53004 10734 53060
rect 15362 53004 15372 53060
rect 15428 53004 22764 53060
rect 22820 53004 22830 53060
rect 27020 52948 27076 53116
rect 31892 53116 33180 53172
rect 33236 53116 33246 53172
rect 41346 53116 41356 53172
rect 41412 53116 42812 53172
rect 42868 53116 42878 53172
rect 31892 53060 31948 53116
rect 29922 53004 29932 53060
rect 29988 53004 31948 53060
rect 32162 53004 32172 53060
rect 32228 53004 36540 53060
rect 36596 53004 36606 53060
rect 9874 52892 9884 52948
rect 9940 52892 10556 52948
rect 10612 52892 11116 52948
rect 11172 52892 11182 52948
rect 23986 52892 23996 52948
rect 24052 52892 25452 52948
rect 25508 52892 26684 52948
rect 26740 52892 26750 52948
rect 27010 52892 27020 52948
rect 27076 52892 27086 52948
rect 30706 52892 30716 52948
rect 30772 52892 31836 52948
rect 31892 52892 31902 52948
rect 33842 52892 33852 52948
rect 33908 52892 37100 52948
rect 37156 52892 37166 52948
rect 1698 52780 1708 52836
rect 1764 52780 2492 52836
rect 2548 52780 2558 52836
rect 18162 52780 18172 52836
rect 18228 52780 19964 52836
rect 20020 52780 20030 52836
rect 35970 52780 35980 52836
rect 36036 52780 40348 52836
rect 40404 52780 41132 52836
rect 41188 52780 41198 52836
rect 42578 52780 42588 52836
rect 42644 52780 44940 52836
rect 44996 52780 45006 52836
rect 10434 52668 10444 52724
rect 10500 52668 11004 52724
rect 11060 52668 11676 52724
rect 11732 52668 11742 52724
rect 12786 52668 12796 52724
rect 12852 52668 14812 52724
rect 14868 52668 15372 52724
rect 15428 52668 24780 52724
rect 24836 52668 24846 52724
rect 19058 52556 19068 52612
rect 19124 52556 26460 52612
rect 26516 52556 26526 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 16706 52444 16716 52500
rect 16772 52444 26908 52500
rect 36306 52444 36316 52500
rect 36372 52444 37324 52500
rect 37380 52444 41244 52500
rect 41300 52444 41310 52500
rect 26852 52388 26908 52444
rect 10210 52332 10220 52388
rect 10276 52332 12460 52388
rect 12516 52332 12526 52388
rect 18284 52332 18396 52388
rect 18452 52332 19068 52388
rect 19124 52332 19134 52388
rect 22092 52332 25228 52388
rect 25284 52332 25294 52388
rect 26852 52332 38668 52388
rect 38724 52332 38734 52388
rect 0 52276 800 52304
rect 0 52220 1708 52276
rect 1764 52220 1774 52276
rect 10322 52220 10332 52276
rect 10388 52220 12796 52276
rect 12852 52220 12862 52276
rect 14578 52220 14588 52276
rect 14644 52220 16492 52276
rect 16548 52220 17276 52276
rect 17332 52220 17948 52276
rect 18004 52220 18014 52276
rect 0 52192 800 52220
rect 18284 52164 18340 52332
rect 22092 52276 22148 52332
rect 20738 52220 20748 52276
rect 20804 52220 21420 52276
rect 21476 52220 22092 52276
rect 22148 52220 22158 52276
rect 23090 52220 23100 52276
rect 23156 52220 27020 52276
rect 27076 52220 27086 52276
rect 31892 52220 32732 52276
rect 32788 52220 32798 52276
rect 36194 52220 36204 52276
rect 36260 52220 36988 52276
rect 37044 52220 37054 52276
rect 31892 52164 31948 52220
rect 11330 52108 11340 52164
rect 11396 52108 12348 52164
rect 12404 52108 18340 52164
rect 25218 52108 25228 52164
rect 25284 52108 29372 52164
rect 29428 52108 29438 52164
rect 29596 52108 31948 52164
rect 34850 52108 34860 52164
rect 34916 52108 35980 52164
rect 36036 52108 36046 52164
rect 37202 52108 37212 52164
rect 37268 52108 38220 52164
rect 38276 52108 38286 52164
rect 29596 52052 29652 52108
rect 23538 51996 23548 52052
rect 23604 51996 25452 52052
rect 25508 51996 26236 52052
rect 26292 51996 26302 52052
rect 26450 51996 26460 52052
rect 26516 51996 26684 52052
rect 26740 51996 29484 52052
rect 29540 51996 29652 52052
rect 39106 51996 39116 52052
rect 39172 51996 42140 52052
rect 42196 51996 42206 52052
rect 3826 51884 3836 51940
rect 3892 51884 10108 51940
rect 10164 51884 10174 51940
rect 15474 51884 15484 51940
rect 15540 51884 16828 51940
rect 16884 51884 18172 51940
rect 18228 51884 18238 51940
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 10882 51660 10892 51716
rect 10948 51660 12068 51716
rect 37314 51660 37324 51716
rect 37380 51660 38108 51716
rect 38164 51660 40180 51716
rect 12012 51604 12068 51660
rect 40124 51604 40180 51660
rect 10770 51548 10780 51604
rect 10836 51548 11564 51604
rect 11620 51548 11630 51604
rect 12002 51548 12012 51604
rect 12068 51548 15036 51604
rect 15092 51548 15102 51604
rect 37986 51548 37996 51604
rect 38052 51548 38892 51604
rect 38948 51548 38958 51604
rect 40114 51548 40124 51604
rect 40180 51548 42252 51604
rect 42308 51548 42318 51604
rect 2034 51436 2044 51492
rect 2100 51436 2716 51492
rect 2772 51436 2782 51492
rect 5618 51436 5628 51492
rect 5684 51436 23548 51492
rect 23604 51436 23614 51492
rect 39666 51436 39676 51492
rect 39732 51436 40908 51492
rect 40964 51436 40974 51492
rect 4386 51324 4396 51380
rect 4452 51324 5180 51380
rect 5236 51324 7644 51380
rect 7700 51324 8988 51380
rect 9044 51324 13132 51380
rect 13188 51324 16604 51380
rect 16660 51324 18732 51380
rect 18788 51324 18798 51380
rect 39442 51324 39452 51380
rect 39508 51324 39518 51380
rect 39452 51268 39508 51324
rect 1810 51212 1820 51268
rect 1876 51212 2492 51268
rect 2548 51212 2558 51268
rect 5058 51212 5068 51268
rect 5124 51212 11900 51268
rect 11956 51212 11966 51268
rect 25890 51212 25900 51268
rect 25956 51212 27580 51268
rect 27636 51212 28252 51268
rect 28308 51212 28318 51268
rect 32610 51212 32620 51268
rect 32676 51212 38556 51268
rect 38612 51212 40348 51268
rect 40404 51212 40414 51268
rect 39218 51100 39228 51156
rect 39284 51100 41468 51156
rect 41524 51100 41534 51156
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 5842 50764 5852 50820
rect 5908 50764 7308 50820
rect 7364 50764 7374 50820
rect 15810 50764 15820 50820
rect 15876 50764 16828 50820
rect 16884 50764 17388 50820
rect 17444 50764 30268 50820
rect 30324 50764 30334 50820
rect 1698 50652 1708 50708
rect 1764 50652 2044 50708
rect 2100 50652 2110 50708
rect 26674 50652 26684 50708
rect 26740 50652 27356 50708
rect 27412 50652 27422 50708
rect 42466 50652 42476 50708
rect 42532 50652 44156 50708
rect 44212 50652 44222 50708
rect 17714 50540 17724 50596
rect 17780 50540 18172 50596
rect 18228 50540 18238 50596
rect 24546 50540 24556 50596
rect 24612 50540 25452 50596
rect 25508 50540 25518 50596
rect 26002 50540 26012 50596
rect 26068 50540 26796 50596
rect 26852 50540 26862 50596
rect 36418 50540 36428 50596
rect 36484 50540 37324 50596
rect 37380 50540 40908 50596
rect 40964 50540 41356 50596
rect 41412 50540 41422 50596
rect 0 50484 800 50512
rect 0 50428 1708 50484
rect 1764 50428 1774 50484
rect 23202 50428 23212 50484
rect 23268 50428 24724 50484
rect 41122 50428 41132 50484
rect 41188 50428 42028 50484
rect 42084 50428 42094 50484
rect 0 50400 800 50428
rect 24668 50372 24724 50428
rect 16006 50316 16044 50372
rect 16100 50316 16110 50372
rect 24658 50316 24668 50372
rect 24724 50316 24734 50372
rect 22754 50204 22764 50260
rect 22820 50204 26236 50260
rect 26292 50204 26302 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 2258 49980 2268 50036
rect 2324 49980 2716 50036
rect 2772 49980 2782 50036
rect 11106 49980 11116 50036
rect 11172 49980 12012 50036
rect 12068 49980 12078 50036
rect 14354 49980 14364 50036
rect 14420 49980 15260 50036
rect 15316 49980 16268 50036
rect 16324 49980 16604 50036
rect 16660 49980 16670 50036
rect 32498 49980 32508 50036
rect 32564 49980 33180 50036
rect 33236 49980 33246 50036
rect 3826 49868 3836 49924
rect 3892 49868 10780 49924
rect 10836 49868 10846 49924
rect 18386 49868 18396 49924
rect 18452 49868 22204 49924
rect 22260 49868 22270 49924
rect 26852 49868 38444 49924
rect 38500 49868 38510 49924
rect 8530 49756 8540 49812
rect 8596 49756 10444 49812
rect 10500 49756 10510 49812
rect 12226 49756 12236 49812
rect 12292 49756 12572 49812
rect 12628 49756 13132 49812
rect 13188 49756 13198 49812
rect 7970 49644 7980 49700
rect 8036 49644 8876 49700
rect 8932 49644 8942 49700
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 10444 49364 10500 49756
rect 26852 49700 26908 49868
rect 15698 49644 15708 49700
rect 15764 49644 21756 49700
rect 21812 49644 25788 49700
rect 25844 49644 26908 49700
rect 13010 49420 13020 49476
rect 13076 49420 24332 49476
rect 24388 49420 24398 49476
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 10444 49308 11228 49364
rect 11284 49308 11294 49364
rect 12450 49308 12460 49364
rect 12516 49308 12908 49364
rect 12964 49308 28588 49364
rect 28644 49308 28654 49364
rect 15026 49196 15036 49252
rect 15092 49196 16492 49252
rect 16548 49196 20524 49252
rect 20580 49196 21532 49252
rect 21588 49196 21598 49252
rect 31892 49196 32844 49252
rect 32900 49196 34188 49252
rect 34244 49196 34254 49252
rect 31892 49140 31948 49196
rect 10546 49084 10556 49140
rect 10612 49084 28140 49140
rect 28196 49084 28206 49140
rect 30594 49084 30604 49140
rect 30660 49084 31948 49140
rect 32050 49084 32060 49140
rect 32116 49084 33068 49140
rect 33124 49084 33134 49140
rect 17490 48972 17500 49028
rect 17556 48972 18284 49028
rect 18340 48972 19068 49028
rect 19124 48972 19134 49028
rect 19954 48972 19964 49028
rect 20020 48972 21868 49028
rect 21924 48972 21934 49028
rect 24658 48972 24668 49028
rect 24724 48972 27132 49028
rect 27188 48972 27198 49028
rect 27906 48972 27916 49028
rect 27972 48972 32340 49028
rect 34290 48972 34300 49028
rect 34356 48972 35084 49028
rect 35140 48972 35150 49028
rect 35410 48972 35420 49028
rect 35476 48972 35980 49028
rect 36036 48972 36046 49028
rect 43652 48972 45388 49028
rect 45444 48972 45454 49028
rect 32284 48916 32340 48972
rect 43652 48916 43708 48972
rect 8194 48860 8204 48916
rect 8260 48860 15372 48916
rect 15428 48860 15438 48916
rect 17826 48860 17836 48916
rect 17892 48860 19628 48916
rect 19684 48860 19694 48916
rect 20402 48860 20412 48916
rect 20468 48860 29260 48916
rect 29316 48860 32060 48916
rect 32116 48860 32126 48916
rect 32284 48860 43708 48916
rect 10322 48748 10332 48804
rect 10388 48748 11004 48804
rect 11060 48748 11070 48804
rect 13580 48748 14364 48804
rect 14420 48748 14430 48804
rect 15810 48748 15820 48804
rect 15876 48748 16156 48804
rect 16212 48748 16222 48804
rect 19628 48748 19740 48804
rect 19796 48748 19806 48804
rect 31826 48748 31836 48804
rect 31892 48748 32956 48804
rect 33012 48748 33022 48804
rect 33282 48748 33292 48804
rect 33348 48748 34636 48804
rect 34692 48748 34702 48804
rect 0 48692 800 48720
rect 0 48636 1708 48692
rect 1764 48636 2492 48692
rect 2548 48636 2558 48692
rect 0 48608 800 48636
rect 13580 48580 13636 48748
rect 16006 48636 16044 48692
rect 16100 48636 16110 48692
rect 19628 48580 19684 48748
rect 27346 48636 27356 48692
rect 27412 48636 27804 48692
rect 27860 48636 28700 48692
rect 28756 48636 28766 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 13570 48524 13580 48580
rect 13636 48524 13646 48580
rect 14018 48524 14028 48580
rect 14084 48524 14420 48580
rect 18498 48524 18508 48580
rect 18564 48524 19684 48580
rect 25330 48524 25340 48580
rect 25396 48524 27468 48580
rect 27524 48524 27534 48580
rect 28018 48524 28028 48580
rect 28084 48524 33068 48580
rect 33124 48524 33134 48580
rect 2706 48412 2716 48468
rect 2772 48412 3052 48468
rect 3108 48412 3500 48468
rect 3556 48412 3566 48468
rect 8306 48412 8316 48468
rect 8372 48412 9660 48468
rect 9716 48412 9726 48468
rect 14364 48356 14420 48524
rect 23202 48412 23212 48468
rect 23268 48412 23884 48468
rect 23940 48412 23950 48468
rect 35634 48412 35644 48468
rect 35700 48412 36316 48468
rect 36372 48412 36382 48468
rect 12114 48300 12124 48356
rect 12180 48300 14364 48356
rect 14420 48300 14430 48356
rect 22418 48300 22428 48356
rect 22484 48300 22988 48356
rect 23044 48300 23054 48356
rect 29810 48300 29820 48356
rect 29876 48300 38892 48356
rect 38948 48300 38958 48356
rect 6626 48188 6636 48244
rect 6692 48188 7084 48244
rect 7140 48188 7150 48244
rect 14466 48188 14476 48244
rect 14532 48188 15148 48244
rect 15204 48188 15932 48244
rect 15988 48188 15998 48244
rect 22082 48188 22092 48244
rect 22148 48188 22158 48244
rect 22306 48188 22316 48244
rect 22372 48188 23436 48244
rect 23492 48188 23996 48244
rect 24052 48188 24556 48244
rect 24612 48188 24622 48244
rect 26562 48188 26572 48244
rect 26628 48188 29036 48244
rect 29092 48188 29102 48244
rect 31490 48188 31500 48244
rect 31556 48188 32172 48244
rect 32228 48188 32238 48244
rect 22092 48132 22148 48188
rect 6066 48076 6076 48132
rect 6132 48076 10668 48132
rect 10724 48076 10734 48132
rect 13346 48076 13356 48132
rect 13412 48076 15260 48132
rect 15316 48076 15326 48132
rect 19842 48076 19852 48132
rect 19908 48076 20524 48132
rect 20580 48076 20590 48132
rect 22092 48076 23884 48132
rect 23940 48076 23950 48132
rect 28578 48076 28588 48132
rect 28644 48076 31724 48132
rect 31780 48076 31790 48132
rect 38210 48076 38220 48132
rect 38276 48076 39676 48132
rect 39732 48076 42812 48132
rect 42868 48076 42878 48132
rect 10668 48020 10724 48076
rect 10668 47964 11340 48020
rect 11396 47964 11406 48020
rect 19394 47964 19404 48020
rect 19460 47964 20300 48020
rect 20356 47964 20366 48020
rect 31602 47964 31612 48020
rect 31668 47964 33516 48020
rect 33572 47964 33582 48020
rect 6402 47852 6412 47908
rect 6468 47852 8204 47908
rect 8260 47852 12684 47908
rect 12740 47852 12750 47908
rect 13122 47852 13132 47908
rect 13188 47852 30268 47908
rect 30324 47852 30334 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 2146 47628 2156 47684
rect 2212 47628 3276 47684
rect 3332 47628 3342 47684
rect 8418 47628 8428 47684
rect 8484 47628 28532 47684
rect 31154 47628 31164 47684
rect 31220 47628 33852 47684
rect 33908 47628 33918 47684
rect 34850 47628 34860 47684
rect 34916 47628 35644 47684
rect 35700 47628 35710 47684
rect 28476 47572 28532 47628
rect 8754 47516 8764 47572
rect 8820 47516 10556 47572
rect 10612 47516 10622 47572
rect 25442 47516 25452 47572
rect 25508 47516 26908 47572
rect 26964 47516 26974 47572
rect 28466 47516 28476 47572
rect 28532 47516 28542 47572
rect 28690 47516 28700 47572
rect 28756 47516 30940 47572
rect 30996 47516 31006 47572
rect 32050 47516 32060 47572
rect 32116 47516 47740 47572
rect 47796 47516 47806 47572
rect 2706 47404 2716 47460
rect 2772 47404 3948 47460
rect 4004 47404 4014 47460
rect 7522 47404 7532 47460
rect 7588 47404 7868 47460
rect 7924 47404 11116 47460
rect 11172 47404 11182 47460
rect 17154 47404 17164 47460
rect 17220 47404 17388 47460
rect 17444 47404 18396 47460
rect 18452 47404 19180 47460
rect 19236 47404 20076 47460
rect 20132 47404 20142 47460
rect 20290 47404 20300 47460
rect 20356 47404 21532 47460
rect 21588 47404 21598 47460
rect 27682 47404 27692 47460
rect 27748 47404 31276 47460
rect 31332 47404 31342 47460
rect 33058 47404 33068 47460
rect 33124 47404 33740 47460
rect 33796 47404 38108 47460
rect 38164 47404 38556 47460
rect 38612 47404 38622 47460
rect 18162 47292 18172 47348
rect 18228 47292 25564 47348
rect 25620 47292 25630 47348
rect 41346 47292 41356 47348
rect 41412 47292 42140 47348
rect 42196 47292 42206 47348
rect 22866 47180 22876 47236
rect 22932 47180 34188 47236
rect 34244 47180 34254 47236
rect 3714 47068 3724 47124
rect 3780 47068 4060 47124
rect 4116 47068 7308 47124
rect 7364 47068 8316 47124
rect 8372 47068 8382 47124
rect 20514 47068 20524 47124
rect 20580 47068 31612 47124
rect 31668 47068 31678 47124
rect 33730 47068 33740 47124
rect 33796 47068 35196 47124
rect 35252 47068 35262 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 10210 46956 10220 47012
rect 10276 46956 11452 47012
rect 11508 46956 11518 47012
rect 15362 46956 15372 47012
rect 15428 46956 16156 47012
rect 16212 46956 16222 47012
rect 21634 46956 21644 47012
rect 21700 46956 22652 47012
rect 22708 46956 22718 47012
rect 27570 46956 27580 47012
rect 27636 46956 30156 47012
rect 30212 46956 32508 47012
rect 32564 46956 33628 47012
rect 33684 46956 33694 47012
rect 38770 46956 38780 47012
rect 38836 46956 39452 47012
rect 39508 46956 39518 47012
rect 0 46900 800 46928
rect 0 46844 1708 46900
rect 1764 46844 2492 46900
rect 2548 46844 2558 46900
rect 4498 46844 4508 46900
rect 4564 46844 9324 46900
rect 9380 46844 10332 46900
rect 10388 46844 10398 46900
rect 14802 46844 14812 46900
rect 14868 46844 14878 46900
rect 30258 46844 30268 46900
rect 30324 46844 34076 46900
rect 34132 46844 34142 46900
rect 0 46816 800 46844
rect 14812 46788 14868 46844
rect 4834 46732 4844 46788
rect 4900 46732 7868 46788
rect 7924 46732 9100 46788
rect 9156 46732 9166 46788
rect 13122 46732 13132 46788
rect 13188 46732 14028 46788
rect 14084 46732 14094 46788
rect 14812 46732 15036 46788
rect 15092 46732 15708 46788
rect 15764 46732 16492 46788
rect 16548 46732 31948 46788
rect 32004 46732 32014 46788
rect 35074 46732 35084 46788
rect 35140 46732 36652 46788
rect 36708 46732 36718 46788
rect 39554 46732 39564 46788
rect 39620 46732 40908 46788
rect 40964 46732 40974 46788
rect 7410 46620 7420 46676
rect 7476 46620 11452 46676
rect 11508 46620 11518 46676
rect 19282 46620 19292 46676
rect 19348 46620 22092 46676
rect 22148 46620 22158 46676
rect 23090 46620 23100 46676
rect 23156 46620 23166 46676
rect 23538 46620 23548 46676
rect 23604 46620 24220 46676
rect 24276 46620 25228 46676
rect 25284 46620 25294 46676
rect 39218 46620 39228 46676
rect 39284 46620 40236 46676
rect 40292 46620 41468 46676
rect 41524 46620 41534 46676
rect 23100 46564 23156 46620
rect 23100 46508 34524 46564
rect 34580 46508 34590 46564
rect 38434 46508 38444 46564
rect 38500 46508 39116 46564
rect 39172 46508 39182 46564
rect 9874 46396 9884 46452
rect 9940 46396 10780 46452
rect 10836 46396 10846 46452
rect 15026 46396 15036 46452
rect 15092 46340 15148 46452
rect 20738 46396 20748 46452
rect 20804 46396 23660 46452
rect 23716 46396 23726 46452
rect 32610 46396 32620 46452
rect 32676 46396 33292 46452
rect 33348 46396 33358 46452
rect 15092 46284 21868 46340
rect 21924 46284 21934 46340
rect 24098 46284 24108 46340
rect 24164 46284 24892 46340
rect 24948 46284 24958 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 10434 46172 10444 46228
rect 10500 46172 10556 46228
rect 10612 46172 10622 46228
rect 14466 46172 14476 46228
rect 14532 46172 15484 46228
rect 15540 46172 22316 46228
rect 22372 46172 22382 46228
rect 26852 46172 30044 46228
rect 30100 46172 30110 46228
rect 26852 46116 26908 46172
rect 7410 46060 7420 46116
rect 7476 46060 26908 46116
rect 29484 46060 32956 46116
rect 33012 46060 33022 46116
rect 9874 45948 9884 46004
rect 9940 45948 11116 46004
rect 11172 45948 11900 46004
rect 11956 45948 11966 46004
rect 16370 45948 16380 46004
rect 16436 45948 17724 46004
rect 17780 45948 20860 46004
rect 20916 45948 20926 46004
rect 29484 45892 29540 46060
rect 32050 45948 32060 46004
rect 32116 45948 50316 46004
rect 50372 45948 50382 46004
rect 8642 45836 8652 45892
rect 8708 45836 9548 45892
rect 9604 45836 10892 45892
rect 10948 45836 10958 45892
rect 17266 45836 17276 45892
rect 17332 45836 18844 45892
rect 18900 45836 18910 45892
rect 20066 45836 20076 45892
rect 20132 45836 21420 45892
rect 21476 45836 22092 45892
rect 22148 45836 22158 45892
rect 22428 45836 29484 45892
rect 29540 45836 29550 45892
rect 31826 45836 31836 45892
rect 31892 45836 38668 45892
rect 38724 45836 38734 45892
rect 22428 45780 22484 45836
rect 4498 45724 4508 45780
rect 4564 45724 9324 45780
rect 9380 45724 9996 45780
rect 10052 45724 10062 45780
rect 10658 45724 10668 45780
rect 10724 45724 11676 45780
rect 11732 45724 11742 45780
rect 17938 45724 17948 45780
rect 18004 45724 21756 45780
rect 21812 45724 21822 45780
rect 22418 45724 22428 45780
rect 22484 45724 22494 45780
rect 24546 45724 24556 45780
rect 24612 45724 27356 45780
rect 27412 45724 27422 45780
rect 33170 45724 33180 45780
rect 33236 45724 34748 45780
rect 34804 45724 34814 45780
rect 7074 45612 7084 45668
rect 7140 45612 8092 45668
rect 8148 45612 8158 45668
rect 15092 45612 28812 45668
rect 28868 45612 28878 45668
rect 32722 45612 32732 45668
rect 32788 45612 34300 45668
rect 34356 45612 34366 45668
rect 35634 45612 35644 45668
rect 35700 45612 38668 45668
rect 38724 45612 39228 45668
rect 39284 45612 39294 45668
rect 6178 45500 6188 45556
rect 6244 45500 6972 45556
rect 7028 45500 7038 45556
rect 10882 45500 10892 45556
rect 10948 45500 11228 45556
rect 11284 45500 11294 45556
rect 15092 45444 15148 45612
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 4162 45388 4172 45444
rect 4228 45388 6524 45444
rect 6580 45388 6748 45444
rect 6804 45388 7980 45444
rect 8036 45388 8046 45444
rect 12002 45388 12012 45444
rect 12068 45388 15148 45444
rect 20738 45388 20748 45444
rect 20804 45388 20972 45444
rect 21028 45388 21038 45444
rect 1698 45276 1708 45332
rect 1764 45276 2492 45332
rect 2548 45276 2558 45332
rect 11190 45276 11228 45332
rect 11284 45276 11294 45332
rect 23314 45276 23324 45332
rect 23380 45276 29372 45332
rect 29428 45276 29438 45332
rect 32162 45276 32172 45332
rect 32228 45276 35644 45332
rect 35700 45276 41020 45332
rect 41076 45276 41086 45332
rect 10210 45164 10220 45220
rect 10276 45164 10668 45220
rect 10724 45164 10734 45220
rect 14802 45164 14812 45220
rect 14868 45164 18956 45220
rect 19012 45164 19516 45220
rect 19572 45164 20748 45220
rect 20804 45164 20814 45220
rect 22978 45164 22988 45220
rect 23044 45164 25900 45220
rect 25956 45164 25966 45220
rect 26338 45164 26348 45220
rect 26404 45164 29148 45220
rect 29204 45164 29214 45220
rect 0 45108 800 45136
rect 0 45052 1708 45108
rect 1764 45052 1774 45108
rect 7746 45052 7756 45108
rect 7812 45052 13692 45108
rect 13748 45052 14364 45108
rect 14420 45052 14430 45108
rect 17266 45052 17276 45108
rect 17332 45052 26124 45108
rect 26180 45052 26190 45108
rect 32498 45052 32508 45108
rect 32564 45052 33404 45108
rect 33460 45052 33470 45108
rect 0 45024 800 45052
rect 3714 44940 3724 44996
rect 3780 44940 8428 44996
rect 8484 44940 8494 44996
rect 9650 44940 9660 44996
rect 9716 44940 10108 44996
rect 10164 44940 10174 44996
rect 10658 44940 10668 44996
rect 10724 44940 11340 44996
rect 11396 44940 11406 44996
rect 19058 44940 19068 44996
rect 19124 44940 20524 44996
rect 20580 44940 20590 44996
rect 23650 44940 23660 44996
rect 23716 44940 24668 44996
rect 24724 44940 25116 44996
rect 25172 44940 25340 44996
rect 25396 44940 25788 44996
rect 25844 44940 25854 44996
rect 41010 44940 41020 44996
rect 41076 44940 44492 44996
rect 44548 44940 44558 44996
rect 10108 44884 10164 44940
rect 1474 44828 1484 44884
rect 1540 44828 3164 44884
rect 3220 44828 3230 44884
rect 10108 44828 15148 44884
rect 18610 44828 18620 44884
rect 18676 44828 20972 44884
rect 21028 44828 21038 44884
rect 15092 44772 15148 44828
rect 6514 44716 6524 44772
rect 6580 44716 7196 44772
rect 7252 44716 10108 44772
rect 10164 44716 10174 44772
rect 15092 44716 15260 44772
rect 15316 44716 15326 44772
rect 19954 44716 19964 44772
rect 20020 44716 22092 44772
rect 22148 44716 23100 44772
rect 23156 44716 23166 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 9762 44604 9772 44660
rect 9828 44604 10220 44660
rect 10276 44604 10286 44660
rect 23986 44604 23996 44660
rect 24052 44604 24444 44660
rect 24500 44604 25116 44660
rect 25172 44604 25182 44660
rect 25778 44604 25788 44660
rect 25844 44604 29820 44660
rect 29876 44604 29886 44660
rect 2230 44492 2268 44548
rect 2324 44492 2334 44548
rect 24668 44492 26908 44548
rect 29922 44492 29932 44548
rect 29988 44492 30940 44548
rect 30996 44492 32396 44548
rect 32452 44492 32462 44548
rect 33842 44492 33852 44548
rect 33908 44492 36204 44548
rect 36260 44492 36270 44548
rect 24668 44436 24724 44492
rect 26852 44436 26908 44492
rect 16930 44380 16940 44436
rect 16996 44380 17612 44436
rect 17668 44380 17678 44436
rect 22194 44380 22204 44436
rect 22260 44380 22652 44436
rect 22708 44380 22718 44436
rect 24658 44380 24668 44436
rect 24724 44380 24734 44436
rect 26852 44380 28140 44436
rect 28196 44380 29148 44436
rect 29204 44380 30380 44436
rect 30436 44380 30446 44436
rect 33506 44380 33516 44436
rect 33572 44380 55356 44436
rect 55412 44380 55422 44436
rect 10098 44268 10108 44324
rect 10164 44268 11004 44324
rect 11060 44268 11070 44324
rect 15698 44268 15708 44324
rect 15764 44268 16380 44324
rect 16436 44268 16446 44324
rect 16818 44268 16828 44324
rect 16884 44268 18060 44324
rect 18116 44268 18126 44324
rect 18386 44268 18396 44324
rect 18452 44268 21420 44324
rect 21476 44268 21486 44324
rect 25218 44268 25228 44324
rect 25284 44268 26236 44324
rect 26292 44268 26302 44324
rect 34738 44268 34748 44324
rect 34804 44268 35420 44324
rect 35476 44268 35486 44324
rect 37090 44268 37100 44324
rect 37156 44268 40012 44324
rect 40068 44268 40908 44324
rect 40964 44268 41580 44324
rect 41636 44268 41646 44324
rect 16380 44212 16436 44268
rect 6850 44156 6860 44212
rect 6916 44156 8092 44212
rect 8148 44156 8158 44212
rect 16380 44156 20300 44212
rect 20356 44156 20366 44212
rect 21858 44156 21868 44212
rect 21924 44156 24780 44212
rect 24836 44156 24846 44212
rect 25078 44156 25116 44212
rect 25172 44156 26572 44212
rect 26628 44156 26638 44212
rect 37426 44156 37436 44212
rect 37492 44156 41020 44212
rect 41076 44156 41086 44212
rect 12786 44044 12796 44100
rect 12852 44044 13692 44100
rect 13748 44044 32060 44100
rect 32116 44044 32126 44100
rect 14018 43932 14028 43988
rect 14084 43932 16604 43988
rect 16660 43932 16670 43988
rect 21410 43932 21420 43988
rect 21476 43932 22092 43988
rect 22148 43932 23436 43988
rect 23492 43932 23502 43988
rect 24322 43932 24332 43988
rect 24388 43932 26572 43988
rect 26628 43932 26638 43988
rect 26852 43932 30604 43988
rect 30660 43932 30670 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 14466 43820 14476 43876
rect 14532 43820 18620 43876
rect 18676 43820 18686 43876
rect 20962 43820 20972 43876
rect 21028 43820 21980 43876
rect 22036 43820 22046 43876
rect 26852 43764 26908 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 8530 43708 8540 43764
rect 8596 43708 11452 43764
rect 11508 43708 11900 43764
rect 11956 43708 12236 43764
rect 12292 43708 12302 43764
rect 16370 43708 16380 43764
rect 16436 43708 17500 43764
rect 17556 43708 17566 43764
rect 18050 43708 18060 43764
rect 18116 43708 19068 43764
rect 19124 43708 19134 43764
rect 22194 43708 22204 43764
rect 22260 43708 26908 43764
rect 33954 43708 33964 43764
rect 34020 43708 37100 43764
rect 37156 43708 37166 43764
rect 39666 43708 39676 43764
rect 39732 43708 41132 43764
rect 41188 43708 41198 43764
rect 1782 43596 1820 43652
rect 1876 43596 1886 43652
rect 3602 43596 3612 43652
rect 3668 43596 4844 43652
rect 4900 43596 5292 43652
rect 5348 43596 6188 43652
rect 6244 43596 6254 43652
rect 7410 43596 7420 43652
rect 7476 43596 11116 43652
rect 11172 43596 12124 43652
rect 12180 43596 12460 43652
rect 12516 43596 12526 43652
rect 17602 43596 17612 43652
rect 17668 43596 18284 43652
rect 18340 43596 19628 43652
rect 19684 43596 19694 43652
rect 26460 43596 29148 43652
rect 29204 43596 29214 43652
rect 31714 43596 31724 43652
rect 31780 43596 31948 43652
rect 33394 43596 33404 43652
rect 33460 43596 34972 43652
rect 35028 43596 35038 43652
rect 37202 43596 37212 43652
rect 37268 43596 38780 43652
rect 38836 43596 39452 43652
rect 39508 43596 39518 43652
rect 40562 43596 40572 43652
rect 40628 43596 41580 43652
rect 41636 43596 41646 43652
rect 26460 43540 26516 43596
rect 2034 43484 2044 43540
rect 2100 43484 2716 43540
rect 2772 43484 2782 43540
rect 7634 43484 7644 43540
rect 7700 43484 8316 43540
rect 8372 43484 8382 43540
rect 9090 43484 9100 43540
rect 9156 43484 13468 43540
rect 13524 43484 13916 43540
rect 13972 43484 13982 43540
rect 15922 43484 15932 43540
rect 15988 43484 18508 43540
rect 18564 43484 18574 43540
rect 21746 43484 21756 43540
rect 21812 43484 22876 43540
rect 22932 43484 24668 43540
rect 24724 43484 26516 43540
rect 26674 43484 26684 43540
rect 26740 43484 27244 43540
rect 27300 43484 27310 43540
rect 30258 43484 30268 43540
rect 30324 43484 30940 43540
rect 30996 43484 31006 43540
rect 31892 43428 31948 43596
rect 40572 43540 40628 43596
rect 33282 43484 33292 43540
rect 33348 43484 37324 43540
rect 37380 43484 37390 43540
rect 39218 43484 39228 43540
rect 39284 43484 40628 43540
rect 5842 43372 5852 43428
rect 5908 43372 6860 43428
rect 6916 43372 7868 43428
rect 7924 43372 7934 43428
rect 8754 43372 8764 43428
rect 8820 43372 10780 43428
rect 10836 43372 10846 43428
rect 12114 43372 12124 43428
rect 12180 43372 12572 43428
rect 12628 43372 12638 43428
rect 15474 43372 15484 43428
rect 15540 43372 17724 43428
rect 17780 43372 17790 43428
rect 25106 43372 25116 43428
rect 25172 43372 26124 43428
rect 26180 43372 26190 43428
rect 26338 43372 26348 43428
rect 26404 43372 28252 43428
rect 28308 43372 28318 43428
rect 31892 43372 32508 43428
rect 32564 43372 33180 43428
rect 33236 43372 33246 43428
rect 0 43316 800 43344
rect 0 43260 1820 43316
rect 1876 43260 1886 43316
rect 33506 43260 33516 43316
rect 33572 43260 38668 43316
rect 38724 43260 38734 43316
rect 0 43232 800 43260
rect 6626 43148 6636 43204
rect 6692 43148 23100 43204
rect 23156 43148 25676 43204
rect 25732 43148 25742 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 24322 43036 24332 43092
rect 24388 43036 24444 43092
rect 24500 43036 24510 43092
rect 24658 42924 24668 42980
rect 24724 42924 27132 42980
rect 27188 42924 27198 42980
rect 33842 42924 33852 42980
rect 33908 42924 44604 42980
rect 44660 42924 44670 42980
rect 10882 42812 10892 42868
rect 10948 42812 20412 42868
rect 20468 42812 20478 42868
rect 21746 42812 21756 42868
rect 21812 42812 22652 42868
rect 22708 42812 22718 42868
rect 33058 42812 33068 42868
rect 33124 42812 34748 42868
rect 34804 42812 35308 42868
rect 35364 42812 35374 42868
rect 8754 42700 8764 42756
rect 8820 42700 10108 42756
rect 10164 42700 10174 42756
rect 11676 42700 17836 42756
rect 17892 42700 17902 42756
rect 22530 42700 22540 42756
rect 22596 42700 22876 42756
rect 22932 42700 22942 42756
rect 23874 42700 23884 42756
rect 23940 42700 24220 42756
rect 24276 42700 24286 42756
rect 28466 42700 28476 42756
rect 28532 42700 29820 42756
rect 29876 42700 30604 42756
rect 30660 42700 30670 42756
rect 35970 42700 35980 42756
rect 36036 42700 36876 42756
rect 36932 42700 40124 42756
rect 40180 42700 40684 42756
rect 40740 42700 40750 42756
rect 11676 42644 11732 42700
rect 2678 42588 2716 42644
rect 2772 42588 2782 42644
rect 8418 42588 8428 42644
rect 8484 42588 9884 42644
rect 9940 42588 9950 42644
rect 10546 42588 10556 42644
rect 10612 42588 11676 42644
rect 11732 42588 11742 42644
rect 12338 42588 12348 42644
rect 12404 42588 27804 42644
rect 27860 42588 27870 42644
rect 3042 42476 3052 42532
rect 3108 42476 3388 42532
rect 7634 42476 7644 42532
rect 7700 42476 11340 42532
rect 11396 42476 11406 42532
rect 18050 42476 18060 42532
rect 18116 42476 21308 42532
rect 21364 42476 21374 42532
rect 3332 42420 3388 42476
rect 3332 42364 18620 42420
rect 18676 42364 18686 42420
rect 26226 42364 26236 42420
rect 26292 42364 30492 42420
rect 30548 42364 30558 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 914 42252 924 42308
rect 980 42252 6300 42308
rect 6356 42252 6366 42308
rect 10210 42252 10220 42308
rect 10276 42252 14028 42308
rect 14084 42252 14094 42308
rect 15092 42252 18060 42308
rect 18116 42252 18126 42308
rect 25340 42252 25452 42308
rect 25508 42252 25518 42308
rect 26338 42252 26348 42308
rect 26404 42252 27020 42308
rect 27076 42252 27086 42308
rect 34514 42252 34524 42308
rect 34580 42252 35420 42308
rect 35476 42252 35486 42308
rect 15092 42196 15148 42252
rect 25340 42196 25396 42252
rect 4050 42140 4060 42196
rect 4116 42140 7308 42196
rect 7364 42140 8652 42196
rect 8708 42140 8718 42196
rect 8866 42140 8876 42196
rect 8932 42140 14364 42196
rect 14420 42140 15148 42196
rect 16706 42140 16716 42196
rect 16772 42140 17612 42196
rect 17668 42140 17678 42196
rect 19394 42140 19404 42196
rect 19460 42140 28588 42196
rect 28644 42140 28654 42196
rect 2230 42028 2268 42084
rect 2324 42028 2334 42084
rect 6402 42028 6412 42084
rect 6468 42028 6972 42084
rect 7028 42028 7644 42084
rect 7700 42028 7710 42084
rect 11778 42028 11788 42084
rect 11844 42028 13916 42084
rect 13972 42028 13982 42084
rect 16594 42028 16604 42084
rect 16660 42028 17948 42084
rect 18004 42028 18014 42084
rect 18498 42028 18508 42084
rect 18564 42028 18844 42084
rect 18900 42028 19964 42084
rect 20020 42028 20748 42084
rect 20804 42028 20814 42084
rect 21074 42028 21084 42084
rect 21140 42028 23100 42084
rect 23156 42028 23166 42084
rect 25890 42028 25900 42084
rect 25956 42028 26348 42084
rect 26404 42028 26414 42084
rect 2034 41916 2044 41972
rect 2100 41916 2716 41972
rect 2772 41916 2782 41972
rect 10406 41916 10444 41972
rect 10500 41916 10510 41972
rect 21970 41916 21980 41972
rect 22036 41916 23436 41972
rect 23492 41916 23502 41972
rect 23986 41916 23996 41972
rect 24052 41916 24556 41972
rect 24612 41916 24622 41972
rect 24770 41916 24780 41972
rect 24836 41916 25676 41972
rect 25732 41916 26236 41972
rect 26292 41916 26302 41972
rect 26562 41916 26572 41972
rect 26628 41916 28700 41972
rect 28756 41916 28766 41972
rect 32050 41916 32060 41972
rect 32116 41916 33964 41972
rect 34020 41916 34524 41972
rect 34580 41916 34590 41972
rect 35522 41916 35532 41972
rect 35588 41916 37772 41972
rect 37828 41916 37838 41972
rect 41346 41916 41356 41972
rect 41412 41916 41422 41972
rect 34524 41860 34580 41916
rect 41356 41860 41412 41916
rect 4050 41804 4060 41860
rect 4116 41804 8652 41860
rect 8708 41804 10556 41860
rect 10612 41804 10622 41860
rect 17826 41804 17836 41860
rect 17892 41804 19852 41860
rect 19908 41804 20300 41860
rect 20356 41804 20366 41860
rect 20962 41804 20972 41860
rect 21028 41804 22484 41860
rect 22866 41804 22876 41860
rect 22932 41804 30940 41860
rect 30996 41804 31006 41860
rect 34524 41804 36316 41860
rect 36372 41804 36382 41860
rect 40114 41804 40124 41860
rect 40180 41804 43820 41860
rect 43876 41804 43886 41860
rect 22428 41748 22484 41804
rect 7522 41692 7532 41748
rect 7588 41692 21532 41748
rect 21588 41692 22204 41748
rect 22260 41692 22270 41748
rect 22428 41692 23100 41748
rect 23156 41692 23166 41748
rect 33842 41692 33852 41748
rect 33908 41692 40012 41748
rect 40068 41692 40078 41748
rect 19506 41580 19516 41636
rect 19572 41580 25788 41636
rect 25844 41580 25854 41636
rect 0 41524 800 41552
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 0 41468 1708 41524
rect 1764 41468 1774 41524
rect 13122 41468 13132 41524
rect 13188 41468 13356 41524
rect 13412 41468 28588 41524
rect 28644 41468 30156 41524
rect 30212 41468 30222 41524
rect 0 41440 800 41468
rect 18834 41356 18844 41412
rect 18900 41356 19628 41412
rect 19684 41356 19694 41412
rect 26226 41356 26236 41412
rect 26292 41356 26908 41412
rect 26964 41356 27580 41412
rect 27636 41356 29372 41412
rect 29428 41356 29438 41412
rect 9538 41244 9548 41300
rect 9604 41244 9996 41300
rect 10052 41244 10062 41300
rect 12450 41244 12460 41300
rect 12516 41244 22876 41300
rect 22932 41244 24332 41300
rect 24388 41244 24780 41300
rect 24836 41244 24846 41300
rect 26852 41244 28140 41300
rect 28196 41244 29148 41300
rect 29204 41244 29214 41300
rect 26852 41188 26908 41244
rect 8082 41132 8092 41188
rect 8148 41132 15148 41188
rect 16370 41132 16380 41188
rect 16436 41132 17612 41188
rect 17668 41132 17678 41188
rect 21382 41132 21420 41188
rect 21476 41132 21486 41188
rect 23202 41132 23212 41188
rect 23268 41132 23996 41188
rect 24052 41132 26908 41188
rect 27570 41132 27580 41188
rect 27636 41132 31388 41188
rect 31444 41132 31454 41188
rect 34626 41132 34636 41188
rect 34692 41132 35420 41188
rect 35476 41132 35486 41188
rect 15092 41076 15148 41132
rect 9650 41020 9660 41076
rect 9716 41020 13692 41076
rect 13748 41020 13758 41076
rect 15092 41020 15708 41076
rect 15764 41020 15774 41076
rect 24770 41020 24780 41076
rect 24836 41020 25900 41076
rect 25956 41020 25966 41076
rect 26786 41020 26796 41076
rect 26852 41020 31164 41076
rect 31220 41020 31230 41076
rect 35186 41020 35196 41076
rect 35252 41020 36876 41076
rect 36932 41020 36942 41076
rect 13906 40908 13916 40964
rect 13972 40908 19852 40964
rect 19908 40908 20524 40964
rect 20580 40908 20590 40964
rect 21074 40908 21084 40964
rect 21140 40908 21980 40964
rect 22036 40908 22046 40964
rect 26674 40908 26684 40964
rect 26740 40908 28476 40964
rect 28532 40908 28542 40964
rect 32946 40908 32956 40964
rect 33012 40908 52668 40964
rect 52724 40908 52734 40964
rect 9538 40796 9548 40852
rect 9604 40796 18172 40852
rect 18228 40796 18620 40852
rect 18676 40796 18686 40852
rect 29362 40796 29372 40852
rect 29428 40796 32172 40852
rect 32228 40796 32238 40852
rect 34514 40796 34524 40852
rect 34580 40796 36204 40852
rect 36260 40796 36270 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 13570 40684 13580 40740
rect 13636 40684 15932 40740
rect 15988 40684 16156 40740
rect 16212 40684 16222 40740
rect 23090 40684 23100 40740
rect 23156 40684 26124 40740
rect 26180 40684 26190 40740
rect 19170 40572 19180 40628
rect 19236 40572 22652 40628
rect 22708 40572 23212 40628
rect 23268 40572 23278 40628
rect 23426 40572 23436 40628
rect 23492 40572 26908 40628
rect 35298 40572 35308 40628
rect 35364 40572 36316 40628
rect 36372 40572 36382 40628
rect 5170 40460 5180 40516
rect 5236 40460 6188 40516
rect 6244 40460 6254 40516
rect 6962 40460 6972 40516
rect 7028 40460 9772 40516
rect 9828 40460 9838 40516
rect 9986 40460 9996 40516
rect 10052 40460 11788 40516
rect 11844 40460 11854 40516
rect 14130 40460 14140 40516
rect 14196 40460 14700 40516
rect 14756 40460 15148 40516
rect 15204 40460 17836 40516
rect 17892 40460 17902 40516
rect 18050 40460 18060 40516
rect 18116 40460 24780 40516
rect 24836 40460 24846 40516
rect 5058 40348 5068 40404
rect 5124 40348 5740 40404
rect 5796 40348 5806 40404
rect 14354 40348 14364 40404
rect 14420 40348 15260 40404
rect 15316 40348 15596 40404
rect 15652 40348 15662 40404
rect 18946 40348 18956 40404
rect 19012 40348 19292 40404
rect 19348 40348 19358 40404
rect 19618 40348 19628 40404
rect 19684 40348 21532 40404
rect 21588 40348 21598 40404
rect 23062 40348 23100 40404
rect 23156 40348 23772 40404
rect 23828 40348 23838 40404
rect 26852 40348 26908 40572
rect 36754 40460 36764 40516
rect 36820 40460 38444 40516
rect 38500 40460 38510 40516
rect 26964 40348 26974 40404
rect 27234 40348 27244 40404
rect 27300 40348 28252 40404
rect 28308 40348 28318 40404
rect 30482 40348 30492 40404
rect 30548 40348 32284 40404
rect 32340 40348 32350 40404
rect 34738 40348 34748 40404
rect 34804 40348 35532 40404
rect 35588 40348 35598 40404
rect 1698 40236 1708 40292
rect 1764 40236 2492 40292
rect 2548 40236 2558 40292
rect 2818 40236 2828 40292
rect 2884 40236 3388 40292
rect 3444 40236 4116 40292
rect 4274 40236 4284 40292
rect 4340 40236 5292 40292
rect 5348 40236 6188 40292
rect 6244 40236 12012 40292
rect 12068 40236 12078 40292
rect 13010 40236 13020 40292
rect 13076 40236 15148 40292
rect 15362 40236 15372 40292
rect 15428 40236 16492 40292
rect 16548 40236 16558 40292
rect 18498 40236 18508 40292
rect 18564 40236 26908 40292
rect 27794 40236 27804 40292
rect 27860 40236 29820 40292
rect 29876 40236 29886 40292
rect 4060 40180 4116 40236
rect 4060 40124 7420 40180
rect 7476 40124 7486 40180
rect 15092 40068 15148 40236
rect 26852 40180 26908 40236
rect 15250 40124 15260 40180
rect 15316 40124 17500 40180
rect 17556 40124 17566 40180
rect 17714 40124 17724 40180
rect 17780 40124 19292 40180
rect 19348 40124 20636 40180
rect 20692 40124 20702 40180
rect 24994 40124 25004 40180
rect 25060 40124 25340 40180
rect 25396 40124 25406 40180
rect 26852 40124 27916 40180
rect 27972 40124 27982 40180
rect 10434 40012 10444 40068
rect 10500 40012 10892 40068
rect 10948 40012 10958 40068
rect 11190 40012 11228 40068
rect 11284 40012 11294 40068
rect 15092 40012 25452 40068
rect 25508 40012 25518 40068
rect 27682 40012 27692 40068
rect 27748 40012 29596 40068
rect 29652 40012 30828 40068
rect 30884 40012 30894 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 4946 39900 4956 39956
rect 5012 39900 6076 39956
rect 6132 39900 28644 39956
rect 28588 39844 28644 39900
rect 2930 39788 2940 39844
rect 2996 39788 4172 39844
rect 4228 39788 4238 39844
rect 19394 39788 19404 39844
rect 19460 39788 24668 39844
rect 24724 39788 24734 39844
rect 25442 39788 25452 39844
rect 25508 39788 25788 39844
rect 25844 39788 25854 39844
rect 26086 39788 26124 39844
rect 26180 39788 26190 39844
rect 28578 39788 28588 39844
rect 28644 39788 28654 39844
rect 30258 39788 30268 39844
rect 30324 39788 30334 39844
rect 0 39732 800 39760
rect 30268 39732 30324 39788
rect 0 39676 1708 39732
rect 1764 39676 1774 39732
rect 8306 39676 8316 39732
rect 8372 39676 15372 39732
rect 15428 39676 15438 39732
rect 17378 39676 17388 39732
rect 17444 39676 30324 39732
rect 0 39648 800 39676
rect 1026 39564 1036 39620
rect 1092 39564 2044 39620
rect 2100 39564 2110 39620
rect 3042 39564 3052 39620
rect 3108 39564 3388 39620
rect 10770 39564 10780 39620
rect 10836 39564 11788 39620
rect 11844 39564 11854 39620
rect 14130 39564 14140 39620
rect 14196 39564 18732 39620
rect 18788 39564 18798 39620
rect 20402 39564 20412 39620
rect 20468 39564 21308 39620
rect 21364 39564 22204 39620
rect 22260 39564 22270 39620
rect 26852 39564 28028 39620
rect 28084 39564 28094 39620
rect 3332 39452 3388 39564
rect 26852 39508 26908 39564
rect 3444 39452 3454 39508
rect 5618 39452 5628 39508
rect 5684 39452 12908 39508
rect 12964 39452 12974 39508
rect 15698 39452 15708 39508
rect 15764 39452 16380 39508
rect 16436 39452 19628 39508
rect 19684 39452 19694 39508
rect 25554 39452 25564 39508
rect 25620 39452 26348 39508
rect 26404 39452 26908 39508
rect 3332 39340 3500 39396
rect 3556 39340 3566 39396
rect 11554 39340 11564 39396
rect 11620 39340 11788 39396
rect 11844 39340 11854 39396
rect 16482 39340 16492 39396
rect 16548 39340 20300 39396
rect 20356 39340 20366 39396
rect 27010 39340 27020 39396
rect 27076 39340 30380 39396
rect 30436 39340 30446 39396
rect 3332 39060 3388 39340
rect 17826 39228 17836 39284
rect 17892 39228 19404 39284
rect 19460 39228 19470 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 3826 39116 3836 39172
rect 3892 39116 4284 39172
rect 4340 39116 4350 39172
rect 4946 39116 4956 39172
rect 5012 39116 7532 39172
rect 7588 39116 7598 39172
rect 19170 39116 19180 39172
rect 19236 39116 19246 39172
rect 21522 39116 21532 39172
rect 21588 39116 22988 39172
rect 23044 39116 23054 39172
rect 19180 39060 19236 39116
rect 2594 39004 2604 39060
rect 2660 39004 3388 39060
rect 3602 39004 3612 39060
rect 3668 39004 5740 39060
rect 5796 39004 5806 39060
rect 8194 39004 8204 39060
rect 8260 39004 11788 39060
rect 11844 39004 11854 39060
rect 13010 39004 13020 39060
rect 13076 39004 13916 39060
rect 13972 39004 13982 39060
rect 14466 39004 14476 39060
rect 14532 39004 18172 39060
rect 18228 39004 18238 39060
rect 19180 39004 21084 39060
rect 21140 39004 21150 39060
rect 21970 39004 21980 39060
rect 22036 39004 26068 39060
rect 31602 39004 31612 39060
rect 31668 39004 31724 39060
rect 31780 39004 31790 39060
rect 35634 39004 35644 39060
rect 35700 39004 36428 39060
rect 36484 39004 36494 39060
rect 3490 38892 3500 38948
rect 3556 38892 5628 38948
rect 5684 38892 5694 38948
rect 7074 38892 7084 38948
rect 7140 38892 7644 38948
rect 7700 38892 7710 38948
rect 13346 38892 13356 38948
rect 13412 38892 20356 38948
rect 3938 38780 3948 38836
rect 4004 38780 5180 38836
rect 5236 38780 5246 38836
rect 6514 38780 6524 38836
rect 6580 38780 10780 38836
rect 10836 38780 10846 38836
rect 11106 38780 11116 38836
rect 11172 38780 15036 38836
rect 15092 38780 15102 38836
rect 19282 38780 19292 38836
rect 19348 38780 19358 38836
rect 5180 38724 5236 38780
rect 5180 38668 6412 38724
rect 6468 38668 7980 38724
rect 8036 38668 8540 38724
rect 8596 38668 8606 38724
rect 12338 38668 12348 38724
rect 12404 38668 15708 38724
rect 15764 38668 16100 38724
rect 18050 38668 18060 38724
rect 18116 38668 18844 38724
rect 18900 38668 18910 38724
rect 4050 38556 4060 38612
rect 4116 38556 14812 38612
rect 14868 38556 14878 38612
rect 14130 38444 14140 38500
rect 14196 38444 14476 38500
rect 14532 38444 14542 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 16044 38388 16100 38668
rect 19292 38612 19348 38780
rect 20300 38724 20356 38892
rect 23492 38892 24220 38948
rect 24276 38892 24286 38948
rect 23492 38836 23548 38892
rect 22418 38780 22428 38836
rect 22484 38780 23324 38836
rect 23380 38780 23548 38836
rect 26012 38836 26068 39004
rect 26226 38892 26236 38948
rect 26292 38892 27468 38948
rect 27524 38892 27534 38948
rect 35746 38892 35756 38948
rect 35812 38892 38220 38948
rect 38276 38892 38286 38948
rect 26012 38780 26908 38836
rect 26964 38780 26974 38836
rect 31938 38780 31948 38836
rect 32004 38780 33628 38836
rect 33684 38780 33694 38836
rect 20300 38668 25564 38724
rect 25620 38668 25630 38724
rect 26562 38668 26572 38724
rect 26628 38668 28252 38724
rect 28308 38668 28318 38724
rect 28476 38668 29036 38724
rect 29092 38668 29102 38724
rect 31154 38668 31164 38724
rect 31220 38668 33852 38724
rect 33908 38668 33918 38724
rect 35522 38668 35532 38724
rect 35588 38668 36988 38724
rect 37044 38668 37436 38724
rect 37492 38668 37502 38724
rect 37762 38668 37772 38724
rect 37828 38668 39900 38724
rect 39956 38668 39966 38724
rect 28476 38612 28532 38668
rect 18358 38556 18396 38612
rect 18452 38556 18462 38612
rect 19282 38556 19292 38612
rect 19348 38556 19358 38612
rect 19730 38556 19740 38612
rect 19796 38556 20300 38612
rect 20356 38556 20366 38612
rect 28102 38556 28140 38612
rect 28196 38556 28532 38612
rect 30482 38556 30492 38612
rect 30548 38556 31052 38612
rect 31108 38556 32508 38612
rect 32564 38556 32956 38612
rect 33012 38556 33516 38612
rect 33572 38556 33582 38612
rect 18498 38444 18508 38500
rect 18564 38444 28028 38500
rect 28084 38444 28094 38500
rect 31378 38444 31388 38500
rect 31444 38444 32396 38500
rect 32452 38444 32462 38500
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 5282 38332 5292 38388
rect 5348 38332 9548 38388
rect 9604 38332 9614 38388
rect 16044 38332 27916 38388
rect 27972 38332 29260 38388
rect 29316 38332 29326 38388
rect 31154 38332 31164 38388
rect 31220 38332 31612 38388
rect 31668 38332 31678 38388
rect 12226 38220 12236 38276
rect 12292 38220 12796 38276
rect 12852 38220 20020 38276
rect 28578 38220 28588 38276
rect 28644 38220 37212 38276
rect 37268 38220 37278 38276
rect 9762 38108 9772 38164
rect 9828 38108 11116 38164
rect 11172 38108 11182 38164
rect 16034 38108 16044 38164
rect 16100 38108 19740 38164
rect 19796 38108 19806 38164
rect 18732 38052 18788 38108
rect 19964 38052 20020 38220
rect 30034 38108 30044 38164
rect 30100 38108 31276 38164
rect 31332 38108 34188 38164
rect 34244 38108 34254 38164
rect 4722 37996 4732 38052
rect 4788 37996 8204 38052
rect 8260 37996 8270 38052
rect 17938 37996 17948 38052
rect 18004 37996 18508 38052
rect 18564 37996 18574 38052
rect 18732 37996 18844 38052
rect 18900 37996 18910 38052
rect 19254 37996 19292 38052
rect 19348 37996 19358 38052
rect 19954 37996 19964 38052
rect 20020 37996 20030 38052
rect 23202 37996 23212 38052
rect 23268 37996 26124 38052
rect 26180 37996 26190 38052
rect 0 37940 800 37968
rect 0 37884 1708 37940
rect 1764 37884 1774 37940
rect 12124 37884 14140 37940
rect 14196 37884 14476 37940
rect 14532 37884 14542 37940
rect 16146 37884 16156 37940
rect 16212 37884 17668 37940
rect 17826 37884 17836 37940
rect 17892 37884 19068 37940
rect 19124 37884 19740 37940
rect 19796 37884 19806 37940
rect 20178 37884 20188 37940
rect 20244 37884 22428 37940
rect 22484 37884 26684 37940
rect 26740 37884 26750 37940
rect 27346 37884 27356 37940
rect 27412 37884 28140 37940
rect 28196 37884 28206 37940
rect 28690 37884 28700 37940
rect 28756 37884 30604 37940
rect 30660 37884 30670 37940
rect 32050 37884 32060 37940
rect 32116 37884 33404 37940
rect 33460 37884 33470 37940
rect 0 37856 800 37884
rect 12124 37828 12180 37884
rect 2006 37772 2044 37828
rect 2100 37772 2110 37828
rect 2790 37772 2828 37828
rect 2884 37772 2894 37828
rect 5618 37772 5628 37828
rect 5684 37772 7084 37828
rect 7140 37772 12124 37828
rect 12180 37772 12190 37828
rect 12338 37772 12348 37828
rect 12404 37772 13692 37828
rect 13748 37772 13758 37828
rect 15810 37772 15820 37828
rect 15876 37772 16828 37828
rect 16884 37772 16894 37828
rect 17612 37716 17668 37884
rect 17938 37772 17948 37828
rect 18004 37772 18172 37828
rect 18228 37772 18238 37828
rect 18946 37772 18956 37828
rect 19012 37772 19628 37828
rect 19684 37772 24108 37828
rect 24164 37772 24174 37828
rect 27570 37772 27580 37828
rect 27636 37772 29708 37828
rect 29764 37772 29774 37828
rect 31714 37772 31724 37828
rect 31780 37772 32172 37828
rect 32228 37772 33292 37828
rect 33348 37772 33852 37828
rect 33908 37772 33918 37828
rect 2370 37660 2380 37716
rect 2436 37660 2716 37716
rect 2772 37660 2782 37716
rect 10658 37660 10668 37716
rect 10724 37660 11116 37716
rect 11172 37660 11182 37716
rect 13010 37660 13020 37716
rect 13076 37660 15036 37716
rect 15092 37660 16548 37716
rect 17612 37660 19684 37716
rect 20850 37660 20860 37716
rect 20916 37660 23436 37716
rect 23492 37660 23502 37716
rect 23874 37660 23884 37716
rect 23940 37660 32116 37716
rect 16492 37604 16548 37660
rect 8978 37548 8988 37604
rect 9044 37548 9212 37604
rect 9268 37548 16156 37604
rect 16212 37548 16222 37604
rect 16482 37548 16492 37604
rect 16548 37548 17500 37604
rect 17556 37548 17566 37604
rect 18284 37548 18508 37604
rect 18564 37548 18574 37604
rect 19366 37548 19404 37604
rect 19460 37548 19470 37604
rect 18284 37492 18340 37548
rect 19628 37492 19684 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 22082 37548 22092 37604
rect 22148 37548 22764 37604
rect 22820 37548 23100 37604
rect 23156 37548 23166 37604
rect 24546 37548 24556 37604
rect 24612 37548 25788 37604
rect 25844 37548 25854 37604
rect 26898 37548 26908 37604
rect 26964 37548 27468 37604
rect 27524 37548 28476 37604
rect 28532 37548 28542 37604
rect 1810 37436 1820 37492
rect 1876 37436 2604 37492
rect 2660 37436 2670 37492
rect 7410 37436 7420 37492
rect 7476 37436 10388 37492
rect 10518 37436 10556 37492
rect 10612 37436 10622 37492
rect 11890 37436 11900 37492
rect 11956 37436 12572 37492
rect 12628 37436 12638 37492
rect 13906 37436 13916 37492
rect 13972 37436 16548 37492
rect 16818 37436 16828 37492
rect 16884 37436 17164 37492
rect 17220 37436 17230 37492
rect 18274 37436 18284 37492
rect 18340 37436 18350 37492
rect 19628 37436 24276 37492
rect 24434 37436 24444 37492
rect 24500 37436 26124 37492
rect 26180 37436 29036 37492
rect 29092 37436 29484 37492
rect 29540 37436 29550 37492
rect 8754 37324 8764 37380
rect 8820 37324 9548 37380
rect 9604 37324 9614 37380
rect 10332 37268 10388 37436
rect 16492 37380 16548 37436
rect 18284 37380 18340 37436
rect 24220 37380 24276 37436
rect 11106 37324 11116 37380
rect 11172 37324 12124 37380
rect 12180 37324 12190 37380
rect 12348 37324 16044 37380
rect 16100 37324 16110 37380
rect 16482 37324 16492 37380
rect 16548 37324 18340 37380
rect 18946 37324 18956 37380
rect 19012 37324 20076 37380
rect 20132 37324 20142 37380
rect 22530 37324 22540 37380
rect 22596 37324 22988 37380
rect 23044 37324 23884 37380
rect 23940 37324 23950 37380
rect 24220 37324 25116 37380
rect 25172 37324 25788 37380
rect 25844 37324 25854 37380
rect 27356 37324 28980 37380
rect 29586 37324 29596 37380
rect 29652 37324 31500 37380
rect 31556 37324 31566 37380
rect 12348 37268 12404 37324
rect 3602 37212 3612 37268
rect 3668 37212 10108 37268
rect 10164 37212 10174 37268
rect 10332 37212 12404 37268
rect 15026 37212 15036 37268
rect 15092 37212 15932 37268
rect 15988 37212 15998 37268
rect 16146 37212 16156 37268
rect 16212 37212 17276 37268
rect 17332 37212 17342 37268
rect 17490 37212 17500 37268
rect 17556 37212 23660 37268
rect 23716 37212 23726 37268
rect 26450 37212 26460 37268
rect 26516 37212 26908 37268
rect 26964 37212 26974 37268
rect 27356 37156 27412 37324
rect 28924 37268 28980 37324
rect 32060 37268 32116 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 32946 37436 32956 37492
rect 33012 37436 38220 37492
rect 38276 37436 39564 37492
rect 39620 37436 39630 37492
rect 28914 37212 28924 37268
rect 28980 37212 29820 37268
rect 29876 37212 29886 37268
rect 32050 37212 32060 37268
rect 32116 37212 32126 37268
rect 32386 37212 32396 37268
rect 32452 37212 34300 37268
rect 34356 37212 36092 37268
rect 36148 37212 36158 37268
rect 1698 37100 1708 37156
rect 1764 37100 3164 37156
rect 3220 37100 3230 37156
rect 3332 37100 17388 37156
rect 17444 37100 17454 37156
rect 19366 37100 19404 37156
rect 19460 37100 19470 37156
rect 20066 37100 20076 37156
rect 20132 37100 22652 37156
rect 22708 37100 22718 37156
rect 23090 37100 23100 37156
rect 23156 37100 27412 37156
rect 27794 37100 27804 37156
rect 27860 37100 28476 37156
rect 28532 37100 29596 37156
rect 29652 37100 29662 37156
rect 30034 37100 30044 37156
rect 30100 37100 31948 37156
rect 32004 37100 32014 37156
rect 3332 37044 3388 37100
rect 2594 36988 2604 37044
rect 2660 36988 3388 37044
rect 11778 36988 11788 37044
rect 11844 36988 13468 37044
rect 13524 36988 13534 37044
rect 15138 36988 15148 37044
rect 15204 36988 16156 37044
rect 16212 36988 16222 37044
rect 16370 36988 16380 37044
rect 16436 36988 16474 37044
rect 16566 36988 16604 37044
rect 16660 36988 16670 37044
rect 20290 36988 20300 37044
rect 20356 36988 22876 37044
rect 22932 36988 22942 37044
rect 25778 36988 25788 37044
rect 25844 36988 30492 37044
rect 30548 36988 30558 37044
rect 15026 36876 15036 36932
rect 15092 36876 18396 36932
rect 18452 36876 19180 36932
rect 19236 36876 19246 36932
rect 21634 36876 21644 36932
rect 21700 36876 23324 36932
rect 23380 36876 23390 36932
rect 36306 36876 36316 36932
rect 36372 36876 36764 36932
rect 36820 36876 36830 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 15474 36764 15484 36820
rect 15540 36764 17164 36820
rect 17220 36764 17230 36820
rect 8642 36652 8652 36708
rect 8708 36652 9996 36708
rect 10052 36652 10062 36708
rect 14130 36652 14140 36708
rect 14196 36652 14924 36708
rect 14980 36652 14990 36708
rect 18050 36652 18060 36708
rect 18116 36652 18620 36708
rect 18676 36652 18686 36708
rect 23874 36652 23884 36708
rect 23940 36652 29148 36708
rect 29204 36652 29214 36708
rect 2006 36540 2044 36596
rect 2100 36540 2110 36596
rect 18834 36540 18844 36596
rect 18900 36540 20748 36596
rect 20804 36540 23996 36596
rect 24052 36540 24062 36596
rect 24210 36540 24220 36596
rect 24276 36540 24314 36596
rect 24406 36540 24444 36596
rect 24500 36540 24510 36596
rect 25890 36540 25900 36596
rect 25956 36540 27580 36596
rect 27636 36540 27646 36596
rect 34626 36540 34636 36596
rect 34692 36540 36092 36596
rect 36148 36540 36652 36596
rect 36708 36540 36718 36596
rect 1586 36428 1596 36484
rect 1652 36428 4620 36484
rect 4676 36428 4686 36484
rect 13122 36428 13132 36484
rect 13188 36428 13804 36484
rect 13860 36428 13870 36484
rect 14354 36428 14364 36484
rect 14420 36428 18060 36484
rect 18116 36428 20860 36484
rect 20916 36428 20926 36484
rect 24098 36428 24108 36484
rect 24164 36428 25452 36484
rect 25508 36428 29708 36484
rect 29764 36428 29774 36484
rect 36306 36428 36316 36484
rect 36372 36428 38892 36484
rect 38948 36428 38958 36484
rect 1932 36372 1988 36428
rect 1922 36316 1932 36372
rect 1988 36316 1998 36372
rect 2930 36316 2940 36372
rect 2996 36316 3276 36372
rect 3332 36316 3836 36372
rect 3892 36316 3902 36372
rect 5954 36316 5964 36372
rect 6020 36316 6748 36372
rect 6804 36316 6814 36372
rect 10210 36316 10220 36372
rect 10276 36316 10444 36372
rect 10500 36316 10892 36372
rect 10948 36316 12572 36372
rect 12628 36316 12638 36372
rect 16594 36316 16604 36372
rect 16660 36316 20188 36372
rect 20244 36316 22876 36372
rect 22932 36316 22942 36372
rect 28018 36316 28028 36372
rect 28084 36316 28364 36372
rect 28420 36316 28430 36372
rect 1362 36204 1372 36260
rect 1428 36204 4284 36260
rect 4340 36204 4844 36260
rect 4900 36204 4910 36260
rect 12114 36204 12124 36260
rect 12180 36204 15148 36260
rect 16258 36204 16268 36260
rect 16324 36204 17836 36260
rect 17892 36204 17902 36260
rect 18508 36204 19740 36260
rect 19796 36204 20412 36260
rect 20468 36204 20478 36260
rect 21298 36204 21308 36260
rect 21364 36204 21980 36260
rect 22036 36204 28476 36260
rect 28532 36204 29260 36260
rect 29316 36204 29326 36260
rect 0 36148 800 36176
rect 0 36092 1708 36148
rect 1764 36092 1774 36148
rect 7980 36092 13580 36148
rect 13636 36092 14980 36148
rect 15092 36092 15148 36204
rect 18508 36148 18564 36204
rect 15204 36092 18564 36148
rect 0 36064 800 36092
rect 7980 36036 8036 36092
rect 14924 36036 14980 36092
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 1922 35980 1932 36036
rect 1988 35980 2716 36036
rect 2772 35980 2782 36036
rect 2930 35980 2940 36036
rect 2996 35980 3276 36036
rect 3332 35980 3342 36036
rect 7970 35980 7980 36036
rect 8036 35980 8046 36036
rect 11330 35980 11340 36036
rect 11396 35980 14196 36036
rect 14924 35980 19404 36036
rect 19460 35980 19470 36036
rect 20636 35980 20748 36036
rect 20804 35980 20814 36036
rect 21522 35980 21532 36036
rect 21588 35980 25620 36036
rect 33506 35980 33516 36036
rect 33572 35980 35532 36036
rect 35588 35980 37660 36036
rect 37716 35980 37726 36036
rect 14140 35924 14196 35980
rect 19404 35924 19460 35980
rect 20636 35924 20692 35980
rect 2594 35868 2604 35924
rect 2660 35868 9996 35924
rect 10052 35868 10062 35924
rect 10406 35868 10444 35924
rect 10500 35868 10668 35924
rect 10724 35868 10734 35924
rect 12002 35868 12012 35924
rect 12068 35868 13916 35924
rect 13972 35868 13982 35924
rect 14140 35868 18396 35924
rect 18452 35868 18462 35924
rect 19404 35868 20692 35924
rect 20850 35868 20860 35924
rect 20916 35868 22876 35924
rect 22932 35868 22942 35924
rect 14802 35756 14812 35812
rect 14868 35756 15148 35812
rect 15250 35756 15260 35812
rect 15316 35756 19012 35812
rect 19170 35756 19180 35812
rect 19236 35756 25340 35812
rect 25396 35756 25406 35812
rect 15092 35700 15148 35756
rect 18956 35700 19012 35756
rect 25564 35700 25620 35980
rect 27010 35868 27020 35924
rect 27076 35868 28700 35924
rect 28756 35868 28766 35924
rect 30146 35868 30156 35924
rect 30212 35868 34748 35924
rect 34804 35868 34814 35924
rect 38098 35868 38108 35924
rect 38164 35868 38668 35924
rect 38724 35868 39340 35924
rect 39396 35868 39406 35924
rect 26898 35756 26908 35812
rect 26964 35756 27580 35812
rect 27636 35756 27646 35812
rect 34850 35756 34860 35812
rect 34916 35756 37324 35812
rect 37380 35756 37772 35812
rect 37828 35756 37838 35812
rect 1138 35644 1148 35700
rect 1204 35644 2716 35700
rect 2772 35644 2782 35700
rect 2930 35644 2940 35700
rect 2996 35644 3276 35700
rect 3332 35644 3342 35700
rect 4050 35644 4060 35700
rect 4116 35644 9660 35700
rect 9716 35644 9726 35700
rect 12114 35644 12124 35700
rect 12180 35644 13020 35700
rect 13076 35644 13086 35700
rect 15092 35644 15428 35700
rect 18956 35644 20412 35700
rect 20468 35644 20478 35700
rect 20626 35644 20636 35700
rect 20692 35644 20972 35700
rect 21028 35644 22540 35700
rect 22596 35644 22606 35700
rect 25564 35644 26908 35700
rect 27766 35644 27804 35700
rect 27860 35644 28252 35700
rect 28308 35644 31724 35700
rect 31780 35644 31790 35700
rect 34066 35644 34076 35700
rect 34132 35644 34142 35700
rect 15372 35588 15428 35644
rect 26852 35588 26908 35644
rect 8978 35532 8988 35588
rect 9044 35532 15148 35588
rect 15204 35532 15214 35588
rect 15362 35532 15372 35588
rect 15428 35532 15438 35588
rect 18386 35532 18396 35588
rect 18452 35532 19852 35588
rect 19908 35532 19918 35588
rect 20748 35532 26684 35588
rect 26740 35532 26750 35588
rect 26852 35532 27132 35588
rect 27188 35532 27198 35588
rect 20748 35476 20804 35532
rect 34076 35476 34132 35644
rect 3826 35420 3836 35476
rect 3892 35420 17724 35476
rect 17780 35420 17790 35476
rect 20738 35420 20748 35476
rect 20804 35420 20814 35476
rect 23426 35420 23436 35476
rect 23492 35420 25788 35476
rect 25844 35420 34132 35476
rect 2818 35308 2828 35364
rect 2884 35308 3052 35364
rect 3108 35308 3118 35364
rect 11554 35308 11564 35364
rect 11620 35308 15148 35364
rect 3266 35252 3276 35308
rect 3332 35252 3370 35308
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 15092 35252 15148 35308
rect 17724 35308 19180 35364
rect 19236 35308 19246 35364
rect 21746 35308 21756 35364
rect 21812 35308 24332 35364
rect 24388 35308 24398 35364
rect 26674 35308 26684 35364
rect 26740 35308 26908 35364
rect 26964 35308 26974 35364
rect 27122 35308 27132 35364
rect 27188 35308 27804 35364
rect 27860 35308 27870 35364
rect 28018 35308 28028 35364
rect 28084 35308 28122 35364
rect 29138 35308 29148 35364
rect 29204 35308 30604 35364
rect 30660 35308 30670 35364
rect 31378 35308 31388 35364
rect 31444 35308 33516 35364
rect 33572 35308 33582 35364
rect 34178 35308 34188 35364
rect 34244 35308 34748 35364
rect 34804 35308 34814 35364
rect 36418 35308 36428 35364
rect 36484 35308 37548 35364
rect 37604 35308 39900 35364
rect 39956 35308 39966 35364
rect 17724 35252 17780 35308
rect 33180 35252 33236 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 2034 35196 2044 35252
rect 2100 35196 2716 35252
rect 2772 35196 2782 35252
rect 6738 35196 6748 35252
rect 6804 35196 7420 35252
rect 7476 35196 8540 35252
rect 8596 35196 8606 35252
rect 9986 35196 9996 35252
rect 10052 35196 10332 35252
rect 10388 35196 14700 35252
rect 14756 35196 14766 35252
rect 15092 35196 16884 35252
rect 17714 35196 17724 35252
rect 17780 35196 17790 35252
rect 20290 35196 20300 35252
rect 20356 35196 21308 35252
rect 21364 35196 21374 35252
rect 23650 35196 23660 35252
rect 23716 35196 30828 35252
rect 30884 35196 30894 35252
rect 33170 35196 33180 35252
rect 33236 35196 33246 35252
rect 16828 35140 16884 35196
rect 6290 35084 6300 35140
rect 6356 35084 11340 35140
rect 11396 35084 12236 35140
rect 12292 35084 12302 35140
rect 13122 35084 13132 35140
rect 13188 35084 13468 35140
rect 13524 35084 13534 35140
rect 16818 35084 16828 35140
rect 16884 35084 16894 35140
rect 18498 35084 18508 35140
rect 18564 35084 23772 35140
rect 23828 35084 25340 35140
rect 25396 35084 25406 35140
rect 28130 35084 28140 35140
rect 28196 35084 29036 35140
rect 29092 35084 29102 35140
rect 2370 34972 2380 35028
rect 2436 34972 2446 35028
rect 5394 34972 5404 35028
rect 5460 34972 8372 35028
rect 9650 34972 9660 35028
rect 9716 34972 13916 35028
rect 13972 34972 17836 35028
rect 17892 34972 19292 35028
rect 19348 34972 19358 35028
rect 22082 34972 22092 35028
rect 22148 34972 23548 35028
rect 23604 34972 23614 35028
rect 26226 34972 26236 35028
rect 26292 34972 27132 35028
rect 27188 34972 27198 35028
rect 2006 34748 2044 34804
rect 2100 34748 2110 34804
rect 2380 34580 2436 34972
rect 8316 34916 8372 34972
rect 6178 34860 6188 34916
rect 6244 34860 7308 34916
rect 7364 34860 8092 34916
rect 8148 34860 8158 34916
rect 8316 34860 11788 34916
rect 11844 34860 11854 34916
rect 12562 34860 12572 34916
rect 12628 34860 13468 34916
rect 13524 34860 13534 34916
rect 16902 34860 16940 34916
rect 16996 34860 17006 34916
rect 19618 34860 19628 34916
rect 19684 34860 19852 34916
rect 19908 34860 19918 34916
rect 20066 34860 20076 34916
rect 20132 34860 20300 34916
rect 20356 34860 20366 34916
rect 20962 34860 20972 34916
rect 21028 34860 28252 34916
rect 28308 34860 28318 34916
rect 30370 34860 30380 34916
rect 30436 34860 31052 34916
rect 31108 34860 31118 34916
rect 32162 34860 32172 34916
rect 32228 34860 33068 34916
rect 33124 34860 35084 34916
rect 35140 34860 35150 34916
rect 11442 34748 11452 34804
rect 11508 34748 13692 34804
rect 13748 34748 13758 34804
rect 14914 34748 14924 34804
rect 14980 34748 15148 34804
rect 15204 34748 15214 34804
rect 18274 34748 18284 34804
rect 18340 34748 18844 34804
rect 18900 34748 22764 34804
rect 22820 34748 22830 34804
rect 23734 34748 23772 34804
rect 23828 34748 24332 34804
rect 24388 34748 26012 34804
rect 26068 34748 29820 34804
rect 29876 34748 29886 34804
rect 30034 34748 30044 34804
rect 30100 34748 30138 34804
rect 31714 34748 31724 34804
rect 31780 34748 37548 34804
rect 37604 34748 37614 34804
rect 2930 34636 2940 34692
rect 2996 34636 3164 34692
rect 3220 34636 5292 34692
rect 5348 34636 5358 34692
rect 17826 34636 17836 34692
rect 17892 34636 18508 34692
rect 18564 34636 18574 34692
rect 19058 34636 19068 34692
rect 19124 34636 19516 34692
rect 19572 34636 22652 34692
rect 22708 34636 22718 34692
rect 22866 34636 22876 34692
rect 22932 34636 26908 34692
rect 27010 34636 27020 34692
rect 27076 34636 27132 34692
rect 27188 34636 27198 34692
rect 27682 34636 27692 34692
rect 27748 34636 28140 34692
rect 28196 34636 29260 34692
rect 29316 34636 29326 34692
rect 30146 34636 30156 34692
rect 30212 34636 30222 34692
rect 30370 34636 30380 34692
rect 30436 34636 30940 34692
rect 30996 34636 34636 34692
rect 34692 34636 34702 34692
rect 26852 34580 26908 34636
rect 2380 34524 2492 34580
rect 2548 34524 2558 34580
rect 9650 34524 9660 34580
rect 9716 34524 10556 34580
rect 10612 34524 10622 34580
rect 15026 34524 15036 34580
rect 15092 34524 18060 34580
rect 18116 34524 18126 34580
rect 20374 34524 20412 34580
rect 20468 34524 23548 34580
rect 23604 34524 23614 34580
rect 26852 34524 28252 34580
rect 28308 34524 28318 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 30156 34468 30212 34636
rect 36306 34524 36316 34580
rect 36372 34524 37436 34580
rect 37492 34524 41916 34580
rect 41972 34524 41982 34580
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 1586 34412 1596 34468
rect 1652 34412 12012 34468
rect 12068 34412 12078 34468
rect 14354 34412 14364 34468
rect 14420 34412 14812 34468
rect 14868 34412 14878 34468
rect 15250 34412 15260 34468
rect 15316 34412 19068 34468
rect 19124 34412 19134 34468
rect 20178 34412 20188 34468
rect 20244 34412 30212 34468
rect 34962 34412 34972 34468
rect 35028 34412 35038 34468
rect 0 34356 800 34384
rect 0 34300 1708 34356
rect 1764 34300 2492 34356
rect 2548 34300 2558 34356
rect 4386 34300 4396 34356
rect 4452 34300 5404 34356
rect 5460 34300 5470 34356
rect 10098 34300 10108 34356
rect 10164 34300 10444 34356
rect 10500 34300 10510 34356
rect 12226 34300 12236 34356
rect 12292 34300 17332 34356
rect 18498 34300 18508 34356
rect 18564 34300 25452 34356
rect 25508 34300 25518 34356
rect 0 34272 800 34300
rect 2034 34188 2044 34244
rect 2100 34188 6412 34244
rect 6468 34188 6478 34244
rect 10546 34188 10556 34244
rect 10612 34188 11172 34244
rect 13122 34188 13132 34244
rect 13188 34188 15484 34244
rect 15540 34188 16604 34244
rect 16660 34188 16670 34244
rect 11116 34020 11172 34188
rect 17276 34132 17332 34300
rect 17490 34188 17500 34244
rect 17556 34188 26236 34244
rect 26292 34188 26908 34244
rect 28018 34188 28028 34244
rect 28084 34188 29372 34244
rect 29428 34188 29438 34244
rect 26852 34132 26908 34188
rect 34972 34132 35028 34412
rect 38210 34300 38220 34356
rect 38276 34300 39228 34356
rect 39284 34300 39294 34356
rect 38612 34188 39340 34244
rect 39396 34188 39788 34244
rect 39844 34188 39854 34244
rect 12226 34076 12236 34132
rect 12292 34076 12460 34132
rect 12516 34076 12526 34132
rect 15250 34076 15260 34132
rect 15316 34076 15820 34132
rect 15876 34076 16716 34132
rect 16772 34076 16782 34132
rect 17276 34076 17892 34132
rect 18050 34076 18060 34132
rect 18116 34076 21196 34132
rect 21252 34076 21262 34132
rect 21410 34076 21420 34132
rect 21476 34076 23996 34132
rect 24052 34076 24062 34132
rect 26852 34076 29540 34132
rect 34402 34076 34412 34132
rect 34468 34076 36652 34132
rect 36708 34076 36718 34132
rect 17836 34020 17892 34076
rect 29484 34020 29540 34076
rect 7410 33964 7420 34020
rect 7476 33964 8204 34020
rect 8260 33964 8270 34020
rect 11106 33964 11116 34020
rect 11172 33964 11182 34020
rect 12002 33964 12012 34020
rect 12068 33964 12684 34020
rect 12740 33964 12750 34020
rect 14690 33964 14700 34020
rect 14756 33964 17612 34020
rect 17668 33964 17678 34020
rect 17836 33964 19124 34020
rect 19282 33964 19292 34020
rect 19348 33964 19516 34020
rect 19572 33964 20972 34020
rect 21028 33964 21038 34020
rect 21196 33964 21644 34020
rect 21700 33964 21710 34020
rect 27234 33964 27244 34020
rect 27300 33964 27804 34020
rect 27860 33964 27870 34020
rect 28242 33964 28252 34020
rect 28308 33964 29260 34020
rect 29316 33964 29326 34020
rect 29474 33964 29484 34020
rect 29540 33964 29932 34020
rect 29988 33964 29998 34020
rect 19068 33908 19124 33964
rect 21196 33908 21252 33964
rect 38612 33908 38668 34188
rect 15922 33852 15932 33908
rect 15988 33852 17780 33908
rect 19068 33852 20748 33908
rect 20804 33852 21252 33908
rect 21410 33852 21420 33908
rect 21476 33852 21756 33908
rect 21812 33852 21822 33908
rect 26338 33852 26348 33908
rect 26404 33852 27580 33908
rect 27636 33852 27646 33908
rect 28690 33852 28700 33908
rect 28756 33852 30492 33908
rect 30548 33852 30558 33908
rect 32498 33852 32508 33908
rect 32564 33852 35868 33908
rect 35924 33852 37100 33908
rect 37156 33852 38668 33908
rect 17724 33796 17780 33852
rect 13010 33740 13020 33796
rect 13076 33740 14028 33796
rect 14084 33740 14094 33796
rect 17724 33740 24668 33796
rect 24724 33740 26572 33796
rect 26628 33740 26638 33796
rect 32386 33740 32396 33796
rect 32452 33740 33068 33796
rect 33124 33740 33134 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 11106 33628 11116 33684
rect 11172 33628 17668 33684
rect 20066 33628 20076 33684
rect 20132 33628 20300 33684
rect 20356 33628 20366 33684
rect 20934 33628 20972 33684
rect 21028 33628 21038 33684
rect 25228 33628 25340 33684
rect 25396 33628 26460 33684
rect 26516 33628 27244 33684
rect 27300 33628 27310 33684
rect 3042 33516 3052 33572
rect 3108 33516 4620 33572
rect 4676 33516 4686 33572
rect 16594 33516 16604 33572
rect 16660 33516 17276 33572
rect 17332 33516 17342 33572
rect 17612 33460 17668 33628
rect 25228 33572 25284 33628
rect 17910 33516 17948 33572
rect 18004 33516 18014 33572
rect 21970 33516 21980 33572
rect 22036 33516 24780 33572
rect 24836 33516 25284 33572
rect 26786 33516 26796 33572
rect 26852 33460 26908 33572
rect 27682 33516 27692 33572
rect 27748 33516 28476 33572
rect 28532 33516 28542 33572
rect 30258 33516 30268 33572
rect 30324 33516 30334 33572
rect 33506 33516 33516 33572
rect 33572 33516 34300 33572
rect 34356 33516 34748 33572
rect 34804 33516 34814 33572
rect 38612 33516 40012 33572
rect 40068 33516 41468 33572
rect 41524 33516 41534 33572
rect 30268 33460 30324 33516
rect 3686 33404 3724 33460
rect 3780 33404 3790 33460
rect 10098 33404 10108 33460
rect 10164 33404 10668 33460
rect 10724 33404 17052 33460
rect 17108 33404 17118 33460
rect 17602 33404 17612 33460
rect 17668 33404 19292 33460
rect 19348 33404 19358 33460
rect 19506 33404 19516 33460
rect 19572 33404 19628 33460
rect 19684 33404 19852 33460
rect 19908 33404 19918 33460
rect 23202 33404 23212 33460
rect 23268 33404 25228 33460
rect 25284 33404 25294 33460
rect 26852 33404 30324 33460
rect 32386 33404 32396 33460
rect 32452 33404 33404 33460
rect 33460 33404 34188 33460
rect 34244 33404 34254 33460
rect 38612 33348 38668 33516
rect 5058 33292 5068 33348
rect 5124 33292 5964 33348
rect 6020 33292 6030 33348
rect 9202 33292 9212 33348
rect 9268 33292 9660 33348
rect 9716 33292 12460 33348
rect 12516 33292 12526 33348
rect 13122 33292 13132 33348
rect 13188 33292 21532 33348
rect 21588 33292 23324 33348
rect 23380 33292 27020 33348
rect 27076 33292 28028 33348
rect 28084 33292 28812 33348
rect 28868 33292 28878 33348
rect 37090 33292 37100 33348
rect 37156 33292 37772 33348
rect 37828 33292 38668 33348
rect 1698 33180 1708 33236
rect 1764 33180 2492 33236
rect 2548 33180 2558 33236
rect 12114 33180 12124 33236
rect 12180 33180 12908 33236
rect 12964 33180 16156 33236
rect 16212 33180 16222 33236
rect 17042 33180 17052 33236
rect 17108 33180 21980 33236
rect 22036 33180 22046 33236
rect 22306 33180 22316 33236
rect 22372 33180 23548 33236
rect 23604 33180 25116 33236
rect 25172 33180 25182 33236
rect 26898 33180 26908 33236
rect 26964 33180 27244 33236
rect 27300 33180 27310 33236
rect 28242 33180 28252 33236
rect 28308 33180 29260 33236
rect 29316 33180 29326 33236
rect 2034 33068 2044 33124
rect 2100 33068 3836 33124
rect 3892 33068 3902 33124
rect 7074 33068 7084 33124
rect 7140 33068 14140 33124
rect 14196 33068 14206 33124
rect 14354 33068 14364 33124
rect 14420 33068 14588 33124
rect 14644 33068 16716 33124
rect 16772 33068 16782 33124
rect 17154 33068 17164 33124
rect 17220 33068 18620 33124
rect 18676 33068 18956 33124
rect 19012 33068 19022 33124
rect 19180 33068 20188 33124
rect 20244 33068 20254 33124
rect 22194 33068 22204 33124
rect 22260 33068 22876 33124
rect 22932 33068 22942 33124
rect 23202 33068 23212 33124
rect 23268 33068 23660 33124
rect 23716 33068 23726 33124
rect 27682 33068 27692 33124
rect 27748 33068 29148 33124
rect 29204 33068 29214 33124
rect 30930 33068 30940 33124
rect 30996 33068 31388 33124
rect 31444 33068 35308 33124
rect 35364 33068 35374 33124
rect 37202 33068 37212 33124
rect 37268 33068 38332 33124
rect 38388 33068 38398 33124
rect 14140 33012 14196 33068
rect 19180 33012 19236 33068
rect 12338 32956 12348 33012
rect 12404 32956 13244 33012
rect 13300 32956 13692 33012
rect 13748 32956 13758 33012
rect 14140 32956 15932 33012
rect 15988 32956 15998 33012
rect 16146 32956 16156 33012
rect 16212 32956 16380 33012
rect 16436 32956 19236 33012
rect 21634 32956 21644 33012
rect 21700 32956 23100 33012
rect 23156 32956 23166 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 1026 32844 1036 32900
rect 1092 32844 7644 32900
rect 7700 32844 7710 32900
rect 8866 32844 8876 32900
rect 8932 32844 9660 32900
rect 9716 32844 9726 32900
rect 12898 32844 12908 32900
rect 12964 32844 17612 32900
rect 17668 32844 17678 32900
rect 17826 32844 17836 32900
rect 17892 32844 18284 32900
rect 18340 32844 18350 32900
rect 20626 32844 20636 32900
rect 20692 32844 21868 32900
rect 21924 32844 21934 32900
rect 25452 32844 27468 32900
rect 27524 32844 27534 32900
rect 25452 32788 25508 32844
rect 2818 32732 2828 32788
rect 2884 32732 3388 32788
rect 7746 32732 7756 32788
rect 7812 32732 14924 32788
rect 14980 32732 22428 32788
rect 22484 32732 24668 32788
rect 24724 32732 25452 32788
rect 25508 32732 25518 32788
rect 0 32564 800 32592
rect 3332 32564 3388 32732
rect 9062 32620 9100 32676
rect 9156 32620 9166 32676
rect 10210 32620 10220 32676
rect 10276 32620 14028 32676
rect 14084 32620 14364 32676
rect 14420 32620 16828 32676
rect 16884 32620 17724 32676
rect 17780 32620 17790 32676
rect 26002 32620 26012 32676
rect 26068 32620 27580 32676
rect 27636 32620 28364 32676
rect 28420 32620 28430 32676
rect 33618 32620 33628 32676
rect 33684 32620 33964 32676
rect 34020 32620 39564 32676
rect 39620 32620 39630 32676
rect 0 32508 1708 32564
rect 1764 32508 1774 32564
rect 3332 32508 3612 32564
rect 3668 32508 3678 32564
rect 4946 32508 4956 32564
rect 5012 32508 7308 32564
rect 7364 32508 7374 32564
rect 9202 32508 9212 32564
rect 9268 32508 9884 32564
rect 9940 32508 9950 32564
rect 10294 32508 10332 32564
rect 10388 32508 10398 32564
rect 10770 32508 10780 32564
rect 10836 32508 15148 32564
rect 18834 32508 18844 32564
rect 18900 32508 19068 32564
rect 19124 32508 21980 32564
rect 22036 32508 22046 32564
rect 22866 32508 22876 32564
rect 22932 32508 25340 32564
rect 25396 32508 25406 32564
rect 0 32480 800 32508
rect 4956 32452 5012 32508
rect 15092 32452 15148 32508
rect 1026 32396 1036 32452
rect 1092 32396 5012 32452
rect 12422 32396 12460 32452
rect 12516 32396 12526 32452
rect 13234 32396 13244 32452
rect 13300 32396 13692 32452
rect 13748 32396 14028 32452
rect 14084 32396 14094 32452
rect 15092 32396 15484 32452
rect 15540 32396 15550 32452
rect 15698 32396 15708 32452
rect 15764 32396 23100 32452
rect 23156 32396 23166 32452
rect 35746 32396 35756 32452
rect 35812 32396 37548 32452
rect 37604 32396 37614 32452
rect 6514 32284 6524 32340
rect 6580 32284 10892 32340
rect 10948 32284 10958 32340
rect 15026 32284 15036 32340
rect 15092 32284 17948 32340
rect 18004 32284 18620 32340
rect 18676 32284 18686 32340
rect 19618 32284 19628 32340
rect 19684 32284 27692 32340
rect 27748 32284 27758 32340
rect 19478 32172 19516 32228
rect 19572 32172 19582 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 8642 32060 8652 32116
rect 8708 32060 17836 32116
rect 17892 32060 20412 32116
rect 20468 32060 20478 32116
rect 21298 32060 21308 32116
rect 21364 32060 21420 32116
rect 21476 32060 21486 32116
rect 5618 31948 5628 32004
rect 5684 31948 7084 32004
rect 7140 31948 7150 32004
rect 12114 31948 12124 32004
rect 12180 31948 13132 32004
rect 13188 31948 13198 32004
rect 13794 31948 13804 32004
rect 13860 31948 14924 32004
rect 14980 31948 15148 32004
rect 15204 31948 15214 32004
rect 16482 31948 16492 32004
rect 16548 31948 18172 32004
rect 18228 31948 19628 32004
rect 19684 31948 19964 32004
rect 20020 31948 21420 32004
rect 21476 31948 21644 32004
rect 21700 31948 21710 32004
rect 23202 31948 23212 32004
rect 23268 31948 25564 32004
rect 25620 31948 25630 32004
rect 2258 31836 2268 31892
rect 2324 31836 3500 31892
rect 3556 31836 3566 31892
rect 5954 31836 5964 31892
rect 6020 31836 6972 31892
rect 7028 31836 7038 31892
rect 9090 31836 9100 31892
rect 9156 31836 9548 31892
rect 9604 31836 13580 31892
rect 13636 31836 13646 31892
rect 18274 31836 18284 31892
rect 18340 31836 26908 31892
rect 32050 31836 32060 31892
rect 32116 31836 32396 31892
rect 32452 31836 32462 31892
rect 33058 31836 33068 31892
rect 33124 31836 38668 31892
rect 3042 31724 3052 31780
rect 3108 31724 3388 31780
rect 15446 31724 15484 31780
rect 15540 31724 15820 31780
rect 15876 31724 15886 31780
rect 18498 31724 18508 31780
rect 18564 31724 20188 31780
rect 20244 31724 21868 31780
rect 21924 31724 22428 31780
rect 22484 31724 22494 31780
rect 22866 31724 22876 31780
rect 22932 31724 23660 31780
rect 23716 31724 23726 31780
rect 3332 31556 3388 31724
rect 8082 31612 8092 31668
rect 8148 31612 11452 31668
rect 11508 31612 11518 31668
rect 13906 31612 13916 31668
rect 13972 31612 14812 31668
rect 14868 31612 14878 31668
rect 18946 31612 18956 31668
rect 19012 31612 20076 31668
rect 20132 31612 20580 31668
rect 20738 31612 20748 31668
rect 20804 31612 22204 31668
rect 22260 31612 22270 31668
rect 20524 31556 20580 31612
rect 23660 31556 23716 31724
rect 26852 31668 26908 31836
rect 38612 31780 38668 31836
rect 34514 31724 34524 31780
rect 34580 31724 36988 31780
rect 37044 31724 37884 31780
rect 37940 31724 37950 31780
rect 38612 31724 39116 31780
rect 39172 31724 39182 31780
rect 26852 31612 28028 31668
rect 28084 31612 28094 31668
rect 36082 31612 36092 31668
rect 36148 31612 37324 31668
rect 37380 31612 37390 31668
rect 3332 31500 3948 31556
rect 4004 31500 5516 31556
rect 5572 31500 5582 31556
rect 9090 31500 9100 31556
rect 9156 31500 9436 31556
rect 9492 31500 9884 31556
rect 9940 31500 9950 31556
rect 14914 31500 14924 31556
rect 14980 31500 17836 31556
rect 17892 31500 17902 31556
rect 18050 31500 18060 31556
rect 18116 31500 20300 31556
rect 20356 31500 20366 31556
rect 20524 31500 23604 31556
rect 23660 31500 29708 31556
rect 29764 31500 29774 31556
rect 30930 31500 30940 31556
rect 30996 31500 37212 31556
rect 37268 31500 37278 31556
rect 23548 31444 23604 31500
rect 8418 31388 8428 31444
rect 8484 31388 10892 31444
rect 10948 31388 16604 31444
rect 16660 31388 16670 31444
rect 17938 31388 17948 31444
rect 18004 31388 18956 31444
rect 19012 31388 19022 31444
rect 21410 31388 21420 31444
rect 21476 31388 21486 31444
rect 23548 31388 24220 31444
rect 24276 31388 26684 31444
rect 26740 31388 28476 31444
rect 28532 31388 28542 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 6066 31276 6076 31332
rect 6132 31276 7420 31332
rect 7476 31276 7486 31332
rect 13346 31276 13356 31332
rect 13412 31276 14140 31332
rect 14196 31276 14812 31332
rect 14868 31276 14878 31332
rect 16706 31276 16716 31332
rect 16772 31276 19628 31332
rect 19684 31276 19694 31332
rect 19628 31220 19684 31276
rect 21420 31220 21476 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 27094 31276 27132 31332
rect 27188 31276 27198 31332
rect 12338 31164 12348 31220
rect 12404 31164 13468 31220
rect 13524 31164 13534 31220
rect 14214 31164 14252 31220
rect 14308 31164 14318 31220
rect 15138 31164 15148 31220
rect 15204 31164 16268 31220
rect 16324 31164 18004 31220
rect 19628 31164 22652 31220
rect 22708 31164 22718 31220
rect 29698 31164 29708 31220
rect 29764 31164 33180 31220
rect 33236 31164 33246 31220
rect 17948 31108 18004 31164
rect 1810 31052 1820 31108
rect 1876 31052 3052 31108
rect 3108 31052 3118 31108
rect 3378 31052 3388 31108
rect 3444 31052 4396 31108
rect 4452 31052 4462 31108
rect 10994 31052 11004 31108
rect 11060 31052 15148 31108
rect 16034 31052 16044 31108
rect 16100 31052 17612 31108
rect 17668 31052 17678 31108
rect 17948 31052 18900 31108
rect 19058 31052 19068 31108
rect 19124 31052 20076 31108
rect 20132 31052 20142 31108
rect 22530 31052 22540 31108
rect 22596 31052 22876 31108
rect 22932 31052 22942 31108
rect 34066 31052 34076 31108
rect 34132 31052 35756 31108
rect 35812 31052 35822 31108
rect 15092 30996 15148 31052
rect 18844 30996 18900 31052
rect 2118 30940 2156 30996
rect 2212 30940 2222 30996
rect 8978 30940 8988 30996
rect 9044 30940 10108 30996
rect 10164 30940 11452 30996
rect 11508 30940 11518 30996
rect 15092 30940 16884 30996
rect 17826 30940 17836 30996
rect 17892 30940 18396 30996
rect 18452 30940 18462 30996
rect 18844 30940 23772 30996
rect 23828 30940 23838 30996
rect 25106 30940 25116 30996
rect 25172 30940 26796 30996
rect 26852 30940 26862 30996
rect 27682 30940 27692 30996
rect 27748 30940 29484 30996
rect 29540 30940 29550 30996
rect 33954 30940 33964 30996
rect 34020 30940 35980 30996
rect 36036 30940 36876 30996
rect 36932 30940 36942 30996
rect 16828 30884 16884 30940
rect 13122 30828 13132 30884
rect 13188 30828 15484 30884
rect 15540 30828 15550 30884
rect 16034 30828 16044 30884
rect 16100 30828 16268 30884
rect 16324 30828 16334 30884
rect 16828 30828 17724 30884
rect 17780 30828 17790 30884
rect 18134 30828 18172 30884
rect 18228 30828 18238 30884
rect 18834 30828 18844 30884
rect 18900 30828 26348 30884
rect 26404 30828 26414 30884
rect 0 30772 800 30800
rect 0 30716 1708 30772
rect 1764 30716 1774 30772
rect 14690 30716 14700 30772
rect 14756 30716 19516 30772
rect 19572 30716 19582 30772
rect 19954 30716 19964 30772
rect 20020 30716 21420 30772
rect 21476 30716 27916 30772
rect 27972 30716 27982 30772
rect 0 30688 800 30716
rect 19180 30660 19236 30716
rect 14802 30604 14812 30660
rect 14868 30604 15484 30660
rect 15540 30604 15550 30660
rect 16818 30604 16828 30660
rect 16884 30604 18956 30660
rect 19012 30604 19022 30660
rect 19180 30604 19292 30660
rect 19348 30604 19358 30660
rect 20850 30604 20860 30660
rect 20916 30604 21868 30660
rect 21924 30604 21934 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 6962 30492 6972 30548
rect 7028 30492 7532 30548
rect 7588 30492 15036 30548
rect 15092 30492 15102 30548
rect 17266 30492 17276 30548
rect 17332 30492 17948 30548
rect 18004 30492 18014 30548
rect 22418 30492 22428 30548
rect 22484 30492 22876 30548
rect 22932 30492 22942 30548
rect 11666 30380 11676 30436
rect 11732 30380 19964 30436
rect 20020 30380 20030 30436
rect 21970 30380 21980 30436
rect 22036 30380 24668 30436
rect 24724 30380 24734 30436
rect 2034 30268 2044 30324
rect 2100 30268 6188 30324
rect 6244 30268 6254 30324
rect 15092 30268 16268 30324
rect 16324 30268 16334 30324
rect 19590 30268 19628 30324
rect 19684 30268 19694 30324
rect 22876 30268 23212 30324
rect 23268 30268 23278 30324
rect 24322 30268 24332 30324
rect 24388 30268 25116 30324
rect 25172 30268 25182 30324
rect 36194 30268 36204 30324
rect 36260 30268 38220 30324
rect 38276 30268 38286 30324
rect 15092 30212 15148 30268
rect 22876 30212 22932 30268
rect 3714 30156 3724 30212
rect 3780 30156 6412 30212
rect 6468 30156 7868 30212
rect 7924 30156 7934 30212
rect 8418 30156 8428 30212
rect 8484 30156 11900 30212
rect 11956 30156 12684 30212
rect 12740 30156 12750 30212
rect 13020 30156 15148 30212
rect 16146 30156 16156 30212
rect 16212 30156 18284 30212
rect 18340 30156 18732 30212
rect 18788 30156 21196 30212
rect 21252 30156 21262 30212
rect 21420 30156 22932 30212
rect 23090 30156 23100 30212
rect 23156 30156 23996 30212
rect 24052 30156 25004 30212
rect 25060 30156 25070 30212
rect 25778 30156 25788 30212
rect 25844 30156 26460 30212
rect 26516 30156 26526 30212
rect 28018 30156 28028 30212
rect 28084 30156 28588 30212
rect 28644 30156 28654 30212
rect 30930 30156 30940 30212
rect 30996 30156 31948 30212
rect 32004 30156 32014 30212
rect 34626 30156 34636 30212
rect 34692 30156 34860 30212
rect 34916 30156 35868 30212
rect 35924 30156 36988 30212
rect 37044 30156 37054 30212
rect 13020 30100 13076 30156
rect 21420 30100 21476 30156
rect 4162 30044 4172 30100
rect 4228 30044 5068 30100
rect 5124 30044 8540 30100
rect 8596 30044 8606 30100
rect 9650 30044 9660 30100
rect 9716 30044 10668 30100
rect 10724 30044 10734 30100
rect 11218 30044 11228 30100
rect 11284 30044 12012 30100
rect 12068 30044 12078 30100
rect 12226 30044 12236 30100
rect 12292 30044 12572 30100
rect 12628 30044 12638 30100
rect 13010 30044 13020 30100
rect 13076 30044 13086 30100
rect 14018 30044 14028 30100
rect 14084 30044 17052 30100
rect 17108 30044 17118 30100
rect 19394 30044 19404 30100
rect 19460 30044 19964 30100
rect 20020 30044 20030 30100
rect 20374 30044 20412 30100
rect 20468 30044 21476 30100
rect 21970 30044 21980 30100
rect 22036 30044 23884 30100
rect 23940 30044 25452 30100
rect 25508 30044 25518 30100
rect 25890 30044 25900 30100
rect 25956 30044 26908 30100
rect 28130 30044 28140 30100
rect 28196 30044 31500 30100
rect 31556 30044 31566 30100
rect 26852 29988 26908 30044
rect 2370 29932 2380 29988
rect 2436 29932 3164 29988
rect 3220 29932 3230 29988
rect 5516 29932 5852 29988
rect 5908 29932 5918 29988
rect 6626 29932 6636 29988
rect 6692 29932 16156 29988
rect 16212 29932 16222 29988
rect 19282 29932 19292 29988
rect 19348 29932 22428 29988
rect 22484 29932 22494 29988
rect 23538 29932 23548 29988
rect 23604 29932 25228 29988
rect 25284 29932 25294 29988
rect 26852 29932 30716 29988
rect 30772 29932 30782 29988
rect 3266 29484 3276 29540
rect 3332 29484 3388 29540
rect 3444 29484 3454 29540
rect 5516 29428 5572 29932
rect 5730 29820 5740 29876
rect 5796 29820 7532 29876
rect 7588 29820 7598 29876
rect 11638 29820 11676 29876
rect 11732 29820 11742 29876
rect 13794 29820 13804 29876
rect 13860 29820 14364 29876
rect 14420 29820 14430 29876
rect 20822 29820 20860 29876
rect 20916 29820 20926 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 8530 29708 8540 29764
rect 8596 29708 12012 29764
rect 12068 29708 14924 29764
rect 14980 29708 14990 29764
rect 23762 29708 23772 29764
rect 23828 29708 24220 29764
rect 24276 29708 24286 29764
rect 8082 29596 8092 29652
rect 8148 29596 14812 29652
rect 14868 29596 14878 29652
rect 15670 29596 15708 29652
rect 15764 29596 15774 29652
rect 17938 29596 17948 29652
rect 18004 29596 18956 29652
rect 19012 29596 19022 29652
rect 19506 29596 19516 29652
rect 19572 29596 19740 29652
rect 19796 29596 19806 29652
rect 20066 29596 20076 29652
rect 20132 29596 21308 29652
rect 21364 29596 21374 29652
rect 22642 29596 22652 29652
rect 22708 29596 23436 29652
rect 23492 29596 27244 29652
rect 27300 29596 27804 29652
rect 27860 29596 30380 29652
rect 30436 29596 30446 29652
rect 6066 29484 6076 29540
rect 6132 29484 6412 29540
rect 6468 29484 6478 29540
rect 8642 29484 8652 29540
rect 8708 29484 9772 29540
rect 9828 29484 9838 29540
rect 12114 29484 12124 29540
rect 12180 29484 13692 29540
rect 13748 29484 13758 29540
rect 18610 29484 18620 29540
rect 18676 29484 20412 29540
rect 20468 29484 20478 29540
rect 23762 29484 23772 29540
rect 23828 29484 27468 29540
rect 27524 29484 27534 29540
rect 27906 29484 27916 29540
rect 27972 29484 28588 29540
rect 28644 29484 28654 29540
rect 4610 29372 4620 29428
rect 4676 29372 6188 29428
rect 6244 29372 6254 29428
rect 9650 29372 9660 29428
rect 9716 29372 10668 29428
rect 10724 29372 10734 29428
rect 10994 29372 11004 29428
rect 11060 29372 11788 29428
rect 11844 29372 13132 29428
rect 13188 29372 13198 29428
rect 13906 29372 13916 29428
rect 13972 29372 14364 29428
rect 14420 29372 14430 29428
rect 14802 29372 14812 29428
rect 14868 29372 20188 29428
rect 20244 29372 20254 29428
rect 21746 29372 21756 29428
rect 21812 29372 22204 29428
rect 22260 29372 26908 29428
rect 28354 29372 28364 29428
rect 28420 29372 29036 29428
rect 29092 29372 29708 29428
rect 29764 29372 29774 29428
rect 18722 29260 18732 29316
rect 18788 29260 19964 29316
rect 20020 29260 20030 29316
rect 20738 29260 20748 29316
rect 20804 29260 23548 29316
rect 23604 29260 23614 29316
rect 26852 29204 26908 29372
rect 9090 29148 9100 29204
rect 9156 29148 11228 29204
rect 11284 29148 12124 29204
rect 12180 29148 14924 29204
rect 14980 29148 14990 29204
rect 16380 29148 24332 29204
rect 24388 29148 24398 29204
rect 26852 29148 31836 29204
rect 31892 29148 31902 29204
rect 16380 29092 16436 29148
rect 10770 29036 10780 29092
rect 10836 29036 12348 29092
rect 12404 29036 12414 29092
rect 13682 29036 13692 29092
rect 13748 29036 16436 29092
rect 16594 29036 16604 29092
rect 16660 29036 17500 29092
rect 17556 29036 17566 29092
rect 19282 29036 19292 29092
rect 19348 29036 26348 29092
rect 26404 29036 26414 29092
rect 28690 29036 28700 29092
rect 28756 29036 29484 29092
rect 29540 29036 29550 29092
rect 0 28980 800 29008
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 0 28924 2380 28980
rect 2436 28924 2446 28980
rect 14242 28924 14252 28980
rect 14308 28924 14476 28980
rect 14532 28924 15260 28980
rect 15316 28924 20860 28980
rect 20916 28924 20926 28980
rect 26226 28924 26236 28980
rect 26292 28924 26908 28980
rect 26964 28924 30492 28980
rect 30548 28924 30558 28980
rect 0 28896 800 28924
rect 2230 28812 2268 28868
rect 2324 28812 2334 28868
rect 8866 28812 8876 28868
rect 8932 28812 10556 28868
rect 10612 28812 17500 28868
rect 17556 28812 17566 28868
rect 18834 28812 18844 28868
rect 18900 28812 19516 28868
rect 19572 28812 26684 28868
rect 26740 28812 27580 28868
rect 27636 28812 27646 28868
rect 28802 28812 28812 28868
rect 28868 28812 28878 28868
rect 28812 28756 28868 28812
rect 914 28700 924 28756
rect 980 28700 7532 28756
rect 7588 28700 7598 28756
rect 12674 28700 12684 28756
rect 12740 28700 13356 28756
rect 13412 28700 15148 28756
rect 15204 28700 20076 28756
rect 20132 28700 20142 28756
rect 20412 28700 23212 28756
rect 23268 28700 23278 28756
rect 24546 28700 24556 28756
rect 24612 28700 29260 28756
rect 29316 28700 29326 28756
rect 2258 28588 2268 28644
rect 2324 28588 3388 28644
rect 3444 28588 3948 28644
rect 4004 28588 5740 28644
rect 5796 28588 5806 28644
rect 14914 28588 14924 28644
rect 14980 28588 18844 28644
rect 18900 28588 19292 28644
rect 19348 28588 19358 28644
rect 20412 28532 20468 28700
rect 22642 28588 22652 28644
rect 22708 28588 23324 28644
rect 23380 28588 23390 28644
rect 25106 28588 25116 28644
rect 25172 28588 26012 28644
rect 26068 28588 26078 28644
rect 27458 28588 27468 28644
rect 27524 28588 28364 28644
rect 28420 28588 28430 28644
rect 28578 28588 28588 28644
rect 28644 28588 29148 28644
rect 29204 28588 29596 28644
rect 29652 28588 29662 28644
rect 25116 28532 25172 28588
rect 2034 28476 2044 28532
rect 2100 28476 3276 28532
rect 3332 28476 3342 28532
rect 5170 28476 5180 28532
rect 5236 28476 7980 28532
rect 8036 28476 8046 28532
rect 10210 28476 10220 28532
rect 10276 28476 20468 28532
rect 23426 28476 23436 28532
rect 23492 28476 25172 28532
rect 27570 28476 27580 28532
rect 27636 28476 28028 28532
rect 28084 28476 28094 28532
rect 2230 28364 2268 28420
rect 2324 28364 2334 28420
rect 2930 28364 2940 28420
rect 2996 28364 3500 28420
rect 3556 28364 3566 28420
rect 10322 28364 10332 28420
rect 10388 28364 10780 28420
rect 10836 28364 10846 28420
rect 10994 28364 11004 28420
rect 11060 28364 11452 28420
rect 11508 28364 11518 28420
rect 14914 28364 14924 28420
rect 14980 28364 16604 28420
rect 16660 28364 16670 28420
rect 17042 28364 17052 28420
rect 17108 28364 18284 28420
rect 18340 28364 18732 28420
rect 18788 28364 18798 28420
rect 24322 28364 24332 28420
rect 24388 28364 25452 28420
rect 25508 28364 25518 28420
rect 1474 28252 1484 28308
rect 1540 28252 4732 28308
rect 4788 28252 5740 28308
rect 5796 28252 5806 28308
rect 15138 28252 15148 28308
rect 15204 28252 16716 28308
rect 16772 28252 17164 28308
rect 17220 28252 17230 28308
rect 21634 28252 21644 28308
rect 21700 28252 31052 28308
rect 31108 28252 31118 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 14130 28140 14140 28196
rect 14196 28140 15036 28196
rect 5506 28028 5516 28084
rect 5572 28028 8764 28084
rect 8820 28028 12236 28084
rect 12292 28028 12302 28084
rect 12562 28028 12572 28084
rect 12628 28028 13132 28084
rect 13188 28028 13692 28084
rect 13748 28028 14700 28084
rect 14756 28028 14766 28084
rect 4162 27916 4172 27972
rect 4228 27916 4956 27972
rect 5012 27916 5628 27972
rect 5684 27916 5694 27972
rect 7746 27916 7756 27972
rect 7812 27916 10444 27972
rect 10500 27916 10510 27972
rect 11442 27916 11452 27972
rect 11508 27916 12012 27972
rect 12068 27916 14308 27972
rect 5282 27804 5292 27860
rect 5348 27804 6972 27860
rect 7028 27804 7038 27860
rect 8082 27804 8092 27860
rect 8148 27804 8428 27860
rect 8484 27804 8494 27860
rect 12086 27804 12124 27860
rect 12180 27804 12190 27860
rect 14252 27748 14308 27916
rect 15092 27860 15148 28196
rect 20178 28140 20188 28196
rect 20244 28140 21532 28196
rect 21588 28140 31164 28196
rect 31220 28140 31230 28196
rect 20188 28084 20244 28140
rect 16258 28028 16268 28084
rect 16324 28028 20244 28084
rect 22978 28028 22988 28084
rect 23044 28028 23772 28084
rect 23828 28028 24220 28084
rect 24276 28028 24286 28084
rect 29922 28028 29932 28084
rect 29988 28028 30828 28084
rect 30884 28028 35644 28084
rect 35700 28028 35710 28084
rect 19618 27916 19628 27972
rect 19684 27916 20636 27972
rect 20692 27916 20702 27972
rect 26674 27916 26684 27972
rect 26740 27916 27356 27972
rect 27412 27916 27422 27972
rect 28242 27916 28252 27972
rect 28308 27916 30268 27972
rect 30324 27916 30334 27972
rect 15092 27804 15484 27860
rect 15540 27804 15550 27860
rect 26450 27804 26460 27860
rect 26516 27804 28140 27860
rect 28196 27804 28206 27860
rect 1698 27692 1708 27748
rect 1764 27692 2492 27748
rect 2548 27692 2558 27748
rect 9090 27692 9100 27748
rect 9156 27692 9996 27748
rect 10052 27692 14028 27748
rect 14084 27692 14094 27748
rect 14252 27692 24668 27748
rect 24724 27692 25676 27748
rect 25732 27692 25742 27748
rect 15810 27580 15820 27636
rect 15876 27580 16716 27636
rect 16772 27580 16782 27636
rect 25890 27580 25900 27636
rect 25956 27580 26684 27636
rect 26740 27580 26750 27636
rect 5058 27468 5068 27524
rect 5124 27468 6412 27524
rect 6468 27468 16828 27524
rect 16884 27468 17388 27524
rect 17444 27468 18620 27524
rect 18676 27468 19404 27524
rect 19460 27468 19470 27524
rect 29250 27468 29260 27524
rect 29316 27468 30044 27524
rect 30100 27468 30110 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 10770 27356 10780 27412
rect 10836 27356 14364 27412
rect 14420 27356 14430 27412
rect 14914 27356 14924 27412
rect 14980 27356 15708 27412
rect 15764 27356 17052 27412
rect 17108 27356 17118 27412
rect 18050 27356 18060 27412
rect 18116 27356 18732 27412
rect 18788 27356 18798 27412
rect 2118 27244 2156 27300
rect 2212 27244 2222 27300
rect 3686 27244 3724 27300
rect 3780 27244 3790 27300
rect 4610 27244 4620 27300
rect 4676 27244 17948 27300
rect 18004 27244 22932 27300
rect 0 27188 800 27216
rect 22876 27188 22932 27244
rect 0 27132 1708 27188
rect 1764 27132 1774 27188
rect 6626 27132 6636 27188
rect 6692 27132 9212 27188
rect 9268 27132 9278 27188
rect 12450 27132 12460 27188
rect 12516 27132 18060 27188
rect 18116 27132 18126 27188
rect 18844 27132 21644 27188
rect 21700 27132 21710 27188
rect 22866 27132 22876 27188
rect 22932 27132 23772 27188
rect 23828 27132 24220 27188
rect 24276 27132 24286 27188
rect 0 27104 800 27132
rect 18844 27076 18900 27132
rect 3938 27020 3948 27076
rect 4004 27020 5180 27076
rect 5236 27020 5246 27076
rect 9090 27020 9100 27076
rect 9156 27020 10556 27076
rect 10612 27020 10622 27076
rect 12338 27020 12348 27076
rect 12404 27020 14476 27076
rect 14532 27020 14924 27076
rect 14980 27020 14990 27076
rect 15138 27020 15148 27076
rect 15204 27020 17332 27076
rect 17490 27020 17500 27076
rect 17556 27020 18844 27076
rect 18900 27020 18910 27076
rect 19954 27020 19964 27076
rect 20020 27020 25228 27076
rect 25284 27020 25900 27076
rect 25956 27020 25966 27076
rect 17276 26964 17332 27020
rect 8082 26908 8092 26964
rect 8148 26908 12124 26964
rect 12180 26908 13580 26964
rect 13636 26908 13646 26964
rect 14354 26908 14364 26964
rect 14420 26908 15372 26964
rect 15428 26908 15438 26964
rect 17276 26908 18396 26964
rect 18452 26908 21420 26964
rect 21476 26908 21486 26964
rect 13580 26852 13636 26908
rect 3490 26796 3500 26852
rect 3556 26796 3724 26852
rect 3780 26796 6748 26852
rect 6804 26796 6814 26852
rect 9314 26796 9324 26852
rect 9380 26796 9548 26852
rect 9604 26796 9614 26852
rect 11750 26796 11788 26852
rect 11844 26796 11854 26852
rect 13580 26796 19292 26852
rect 19348 26796 20412 26852
rect 20468 26796 20478 26852
rect 21970 26796 21980 26852
rect 22036 26796 22204 26852
rect 22260 26796 22270 26852
rect 12786 26684 12796 26740
rect 12852 26684 15596 26740
rect 15652 26684 15662 26740
rect 15922 26684 15932 26740
rect 15988 26684 17612 26740
rect 17668 26684 17678 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 9762 26572 9772 26628
rect 9828 26572 10556 26628
rect 10612 26572 10622 26628
rect 14242 26572 14252 26628
rect 14308 26572 19516 26628
rect 19572 26572 19582 26628
rect 25218 26572 25228 26628
rect 25284 26572 27020 26628
rect 27076 26572 27086 26628
rect 5954 26460 5964 26516
rect 6020 26460 9660 26516
rect 9716 26460 9726 26516
rect 10098 26460 10108 26516
rect 10164 26460 11004 26516
rect 11060 26460 11070 26516
rect 12786 26460 12796 26516
rect 12852 26460 13244 26516
rect 13300 26460 13692 26516
rect 13748 26460 13758 26516
rect 15474 26460 15484 26516
rect 15540 26460 21196 26516
rect 21252 26460 21262 26516
rect 21410 26460 21420 26516
rect 21476 26460 26908 26516
rect 15484 26404 15540 26460
rect 26852 26404 26908 26460
rect 5842 26348 5852 26404
rect 5908 26348 7644 26404
rect 7700 26348 7710 26404
rect 10322 26348 10332 26404
rect 10388 26348 15036 26404
rect 15092 26348 15540 26404
rect 15698 26348 15708 26404
rect 15764 26348 16492 26404
rect 16548 26348 16558 26404
rect 17602 26348 17612 26404
rect 17668 26348 18564 26404
rect 20850 26348 20860 26404
rect 20916 26348 25340 26404
rect 25396 26348 25406 26404
rect 26852 26348 27804 26404
rect 27860 26348 28252 26404
rect 28308 26348 28318 26404
rect 18508 26292 18564 26348
rect 9650 26236 9660 26292
rect 9716 26236 11900 26292
rect 11956 26236 13580 26292
rect 13636 26236 13646 26292
rect 16034 26236 16044 26292
rect 16100 26236 17948 26292
rect 18004 26236 18014 26292
rect 18498 26236 18508 26292
rect 18564 26236 25228 26292
rect 25284 26236 25294 26292
rect 10546 26124 10556 26180
rect 10612 26124 16156 26180
rect 16212 26124 16604 26180
rect 16660 26124 17388 26180
rect 17444 26124 17454 26180
rect 22194 26124 22204 26180
rect 22260 26124 23212 26180
rect 23268 26124 23278 26180
rect 5058 26012 5068 26068
rect 5124 26012 5964 26068
rect 6020 26012 6030 26068
rect 7746 26012 7756 26068
rect 7812 26012 10220 26068
rect 10276 26012 10286 26068
rect 10994 26012 11004 26068
rect 11060 26012 15932 26068
rect 15988 26012 15998 26068
rect 16930 26012 16940 26068
rect 16996 26012 19628 26068
rect 19684 26012 19964 26068
rect 20020 26012 23660 26068
rect 23716 26012 23726 26068
rect 20402 25900 20412 25956
rect 20468 25900 25228 25956
rect 25284 25900 25294 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 23090 25788 23100 25844
rect 23156 25788 24220 25844
rect 24276 25788 24286 25844
rect 9538 25676 9548 25732
rect 9604 25676 14084 25732
rect 7298 25564 7308 25620
rect 7364 25564 9660 25620
rect 9716 25564 9726 25620
rect 14028 25508 14084 25676
rect 15260 25676 21420 25732
rect 21476 25676 21486 25732
rect 23426 25676 23436 25732
rect 23492 25676 24444 25732
rect 24500 25676 24510 25732
rect 15260 25620 15316 25676
rect 23436 25620 23492 25676
rect 14914 25564 14924 25620
rect 14980 25564 15260 25620
rect 15316 25564 15326 25620
rect 15810 25564 15820 25620
rect 15876 25564 16380 25620
rect 16436 25564 23492 25620
rect 25218 25564 25228 25620
rect 25284 25564 27132 25620
rect 27188 25564 34860 25620
rect 34916 25564 34926 25620
rect 9090 25452 9100 25508
rect 9156 25452 9436 25508
rect 9492 25452 9502 25508
rect 10994 25452 11004 25508
rect 11060 25452 11900 25508
rect 11956 25452 11966 25508
rect 14018 25452 14028 25508
rect 14084 25452 16044 25508
rect 16100 25452 16716 25508
rect 16772 25452 16782 25508
rect 18498 25452 18508 25508
rect 18564 25452 20972 25508
rect 21028 25452 21038 25508
rect 27906 25452 27916 25508
rect 27972 25452 29260 25508
rect 29316 25452 29326 25508
rect 0 25396 800 25424
rect 0 25340 1708 25396
rect 1764 25340 2492 25396
rect 2548 25340 2558 25396
rect 9538 25340 9548 25396
rect 9604 25340 10444 25396
rect 10500 25340 10510 25396
rect 10770 25340 10780 25396
rect 10836 25340 12572 25396
rect 12628 25340 12638 25396
rect 16818 25340 16828 25396
rect 16884 25340 18844 25396
rect 18900 25340 18910 25396
rect 22754 25340 22764 25396
rect 22820 25340 23548 25396
rect 23604 25340 23614 25396
rect 0 25312 800 25340
rect 11218 25228 11228 25284
rect 11284 25228 12012 25284
rect 12068 25228 13692 25284
rect 13748 25228 15260 25284
rect 15316 25228 15326 25284
rect 17714 25228 17724 25284
rect 17780 25228 18620 25284
rect 18676 25228 18686 25284
rect 19030 25228 19068 25284
rect 19124 25228 20076 25284
rect 20132 25228 21532 25284
rect 21588 25228 22652 25284
rect 22708 25228 22718 25284
rect 13346 25116 13356 25172
rect 13412 25116 13804 25172
rect 13860 25116 13870 25172
rect 17602 25116 17612 25172
rect 17668 25116 17948 25172
rect 18004 25116 18014 25172
rect 23202 25116 23212 25172
rect 23268 25116 24444 25172
rect 24500 25116 24510 25172
rect 26852 25116 29372 25172
rect 29428 25116 29438 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 14018 25004 14028 25060
rect 14084 25004 17388 25060
rect 17444 25004 17454 25060
rect 11666 24892 11676 24948
rect 11732 24892 12348 24948
rect 12404 24892 12414 24948
rect 13010 24892 13020 24948
rect 13076 24892 14700 24948
rect 14756 24892 23772 24948
rect 23828 24892 23838 24948
rect 8754 24780 8764 24836
rect 8820 24780 16940 24836
rect 16996 24780 17006 24836
rect 17154 24780 17164 24836
rect 17220 24780 20244 24836
rect 20850 24780 20860 24836
rect 20916 24780 20972 24836
rect 21028 24780 21532 24836
rect 21588 24780 21598 24836
rect 23314 24780 23324 24836
rect 23380 24780 24220 24836
rect 24276 24780 25004 24836
rect 25060 24780 25070 24836
rect 20188 24724 20244 24780
rect 26852 24724 26908 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 13122 24668 13132 24724
rect 13188 24668 13916 24724
rect 13972 24668 13982 24724
rect 16706 24668 16716 24724
rect 16772 24668 17836 24724
rect 17892 24668 19964 24724
rect 20020 24668 20030 24724
rect 20188 24668 26908 24724
rect 11666 24556 11676 24612
rect 11732 24556 16492 24612
rect 16548 24556 16828 24612
rect 16884 24556 16894 24612
rect 25778 24556 25788 24612
rect 25844 24556 26236 24612
rect 26292 24556 39004 24612
rect 39060 24556 39070 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 15586 24220 15596 24276
rect 15652 24220 16828 24276
rect 16884 24220 27916 24276
rect 27972 24220 27982 24276
rect 15148 24108 21980 24164
rect 22036 24108 22316 24164
rect 22372 24108 22540 24164
rect 22596 24108 22606 24164
rect 15148 24052 15204 24108
rect 9874 23996 9884 24052
rect 9940 23996 15148 24052
rect 15204 23996 15214 24052
rect 19730 23996 19740 24052
rect 19796 23996 21532 24052
rect 21588 23996 21598 24052
rect 24434 23996 24444 24052
rect 24500 23996 25788 24052
rect 25844 23996 25854 24052
rect 20178 23884 20188 23940
rect 20244 23884 21084 23940
rect 21140 23884 21150 23940
rect 24770 23884 24780 23940
rect 24836 23884 25452 23940
rect 25508 23884 25518 23940
rect 2006 23772 2044 23828
rect 2100 23772 2110 23828
rect 12450 23772 12460 23828
rect 12516 23772 15148 23828
rect 15204 23772 15932 23828
rect 15988 23772 15998 23828
rect 16482 23772 16492 23828
rect 16548 23772 18172 23828
rect 18228 23772 18238 23828
rect 19058 23772 19068 23828
rect 19124 23772 24556 23828
rect 24612 23772 25228 23828
rect 25284 23772 25294 23828
rect 0 23604 800 23632
rect 16492 23604 16548 23772
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 11330 23548 11340 23604
rect 11396 23548 16548 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 1138 23436 1148 23492
rect 1204 23436 1820 23492
rect 1876 23436 1886 23492
rect 13346 23436 13356 23492
rect 13412 23436 15148 23492
rect 22418 23436 22428 23492
rect 22484 23436 22494 23492
rect 15092 23380 15148 23436
rect 22428 23380 22484 23436
rect 15092 23324 22484 23380
rect 8306 23212 8316 23268
rect 8372 23044 8428 23268
rect 15810 23212 15820 23268
rect 15876 23212 21308 23268
rect 21364 23212 21374 23268
rect 22194 23212 22204 23268
rect 22260 23212 22988 23268
rect 23044 23212 23054 23268
rect 8372 22988 19068 23044
rect 19124 22988 19134 23044
rect 16146 22876 16156 22932
rect 16212 22876 17612 22932
rect 17668 22876 28028 22932
rect 28084 22876 28094 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 0 21812 800 21840
rect 0 21756 1708 21812
rect 1764 21756 2492 21812
rect 2548 21756 2558 21812
rect 6290 21756 6300 21812
rect 6356 21756 28140 21812
rect 28196 21756 28206 21812
rect 0 21728 800 21756
rect 12226 21644 12236 21700
rect 12292 21644 27804 21700
rect 27860 21644 27870 21700
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 0 20020 800 20048
rect 0 19964 1708 20020
rect 1764 19964 2492 20020
rect 2548 19964 2558 20020
rect 0 19936 800 19964
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 0 18228 800 18256
rect 0 18172 1708 18228
rect 1764 18172 2492 18228
rect 2548 18172 2558 18228
rect 0 18144 800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 0 16436 800 16464
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16380 1708 16436
rect 1764 16380 2492 16436
rect 2548 16380 2558 16436
rect 0 16352 800 16380
rect 1362 15708 1372 15764
rect 1428 15708 1820 15764
rect 1876 15708 1886 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 0 14644 800 14672
rect 0 14588 1708 14644
rect 1764 14588 2492 14644
rect 2548 14588 2558 14644
rect 0 14560 800 14588
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 2034 13356 2044 13412
rect 2100 13356 3836 13412
rect 3892 13356 3902 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 0 12852 800 12880
rect 0 12796 1708 12852
rect 1764 12796 2492 12852
rect 2548 12796 2558 12852
rect 0 12768 800 12796
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 0 11060 800 11088
rect 0 11004 1708 11060
rect 1764 11004 2492 11060
rect 2548 11004 2558 11060
rect 0 10976 800 11004
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 2034 9660 2044 9716
rect 2100 9660 6748 9716
rect 6804 9660 6814 9716
rect 2034 9436 2044 9492
rect 2100 9436 5628 9492
rect 5684 9436 5694 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 0 9268 800 9296
rect 0 9212 1708 9268
rect 1764 9212 2492 9268
rect 2548 9212 2558 9268
rect 0 9184 800 9212
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 1698 7980 1708 8036
rect 1764 7980 2492 8036
rect 2548 7980 2558 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 0 7476 800 7504
rect 0 7420 1708 7476
rect 1764 7420 1774 7476
rect 0 7392 800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 2370 6748 2380 6804
rect 2436 6748 5068 6804
rect 5124 6748 5134 6804
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 1026 5852 1036 5908
rect 1092 5852 2156 5908
rect 2212 5852 2222 5908
rect 0 5684 800 5712
rect 0 5628 1708 5684
rect 1764 5628 1774 5684
rect 0 5600 800 5628
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 0 3892 800 3920
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 0 3836 1708 3892
rect 1764 3836 2492 3892
rect 2548 3836 2558 3892
rect 0 3808 800 3836
rect 1698 3276 1708 3332
rect 1764 3276 2716 3332
rect 2772 3276 2782 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 0 2100 800 2128
rect 0 2044 1708 2100
rect 1764 2044 1774 2100
rect 0 2016 800 2044
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 16044 50316 16100 50372
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 16044 48636 16100 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 10556 46172 10612 46228
rect 15484 46172 15540 46228
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 20972 45388 21028 45444
rect 11228 45276 11284 45332
rect 25116 44940 25172 44996
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 2268 44492 2324 44548
rect 16940 44380 16996 44436
rect 16380 44268 16436 44324
rect 18060 44268 18116 44324
rect 25116 44156 25172 44212
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 1820 43596 1876 43652
rect 12124 43372 12180 43428
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 24444 43036 24500 43092
rect 24220 42700 24276 42756
rect 2716 42588 2772 42644
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 2268 42028 2324 42084
rect 21084 42028 21140 42084
rect 10444 41916 10500 41972
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 12460 41244 12516 41300
rect 21420 41132 21476 41188
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 15932 40684 15988 40740
rect 26124 40684 26180 40740
rect 19180 40572 19236 40628
rect 23100 40348 23156 40404
rect 11228 40012 11284 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 26124 39788 26180 39844
rect 11788 39340 11844 39396
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 21532 39116 21588 39172
rect 18172 39004 18228 39060
rect 31612 39004 31668 39060
rect 15708 38668 15764 38724
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 18396 38556 18452 38612
rect 19292 38556 19348 38612
rect 28140 38556 28196 38612
rect 18508 38444 18564 38500
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 31612 38332 31668 38388
rect 19292 37996 19348 38052
rect 2044 37772 2100 37828
rect 2828 37772 2884 37828
rect 16828 37772 16884 37828
rect 18172 37772 18228 37828
rect 2716 37660 2772 37716
rect 18508 37548 18564 37604
rect 19404 37548 19460 37604
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 1820 37436 1876 37492
rect 10556 37436 10612 37492
rect 25116 37324 25172 37380
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 19404 37100 19460 37156
rect 16380 36988 16436 37044
rect 16604 36988 16660 37044
rect 22876 36988 22932 37044
rect 15036 36876 15092 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 2044 36540 2100 36596
rect 24220 36540 24276 36596
rect 24444 36540 24500 36596
rect 3276 36316 3332 36372
rect 16268 36204 16324 36260
rect 15148 36092 15204 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 10444 35868 10500 35924
rect 20412 35644 20468 35700
rect 27804 35644 27860 35700
rect 2828 35308 2884 35364
rect 3276 35252 3332 35308
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 19180 35308 19236 35364
rect 28028 35308 28084 35364
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 10332 35196 10388 35252
rect 2044 34748 2100 34804
rect 16940 34860 16996 34916
rect 19628 34860 19684 34916
rect 20300 34860 20356 34916
rect 23772 34748 23828 34804
rect 30044 34748 30100 34804
rect 22876 34636 22932 34692
rect 27132 34636 27188 34692
rect 20412 34524 20468 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 20188 34412 20244 34468
rect 12236 34076 12292 34132
rect 21420 33852 21476 33908
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 20300 33628 20356 33684
rect 20972 33628 21028 33684
rect 16604 33516 16660 33572
rect 17948 33516 18004 33572
rect 3724 33404 3780 33460
rect 19628 33404 19684 33460
rect 12460 33292 12516 33348
rect 16716 33068 16772 33124
rect 20188 33068 20244 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 9100 32620 9156 32676
rect 10332 32508 10388 32564
rect 12460 32396 12516 32452
rect 23100 32396 23156 32452
rect 19516 32172 19572 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 21420 32060 21476 32116
rect 19628 31948 19684 32004
rect 15484 31724 15540 31780
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 16716 31276 16772 31332
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 27132 31276 27188 31332
rect 14252 31164 14308 31220
rect 2156 30940 2212 30996
rect 18396 30940 18452 30996
rect 18172 30828 18228 30884
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 15036 30492 15092 30548
rect 11676 30380 11732 30436
rect 16268 30268 16324 30324
rect 19628 30268 19684 30324
rect 20412 30044 20468 30100
rect 11676 29820 11732 29876
rect 20860 29820 20916 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 15708 29596 15764 29652
rect 17948 29596 18004 29652
rect 20412 29484 20468 29540
rect 14924 29148 14980 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 14252 28924 14308 28980
rect 20860 28924 20916 28980
rect 2268 28812 2324 28868
rect 18844 28812 18900 28868
rect 19516 28812 19572 28868
rect 15148 28700 15204 28756
rect 14924 28588 14980 28644
rect 28028 28476 28084 28532
rect 2268 28364 2324 28420
rect 10332 28364 10388 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 15036 28140 15092 28196
rect 12124 27804 12180 27860
rect 23772 28028 23828 28084
rect 30044 27468 30100 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 2156 27244 2212 27300
rect 3724 27244 3780 27300
rect 11788 26796 11844 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 21420 26460 21476 26516
rect 19628 26012 19684 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 21420 25676 21476 25732
rect 9100 25452 9156 25508
rect 20972 25452 21028 25508
rect 18844 25340 18900 25396
rect 19068 25228 19124 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 20860 24780 20916 24836
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 16828 24220 16884 24276
rect 21532 23996 21588 24052
rect 2044 23772 2100 23828
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 19068 22988 19124 23044
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 28140 21756 28196 21812
rect 12236 21644 12292 21700
rect 27804 21644 27860 21700
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 16044 50372 16100 50382
rect 16044 48692 16100 50316
rect 16044 48626 16100 48636
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 2268 44548 2324 44558
rect 1820 43652 1876 43662
rect 1820 37492 1876 43596
rect 2268 42084 2324 44492
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 2268 42018 2324 42028
rect 2716 42644 2772 42654
rect 1820 37426 1876 37436
rect 2044 37828 2100 37838
rect 2044 36596 2100 37772
rect 2716 37716 2772 42588
rect 4448 41580 4768 43092
rect 10556 46228 10612 46238
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 2716 37650 2772 37660
rect 2828 37828 2884 37838
rect 2044 36530 2100 36540
rect 2828 35364 2884 37772
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 2828 35298 2884 35308
rect 3276 36372 3332 36382
rect 3276 35308 3332 36316
rect 3276 35242 3332 35252
rect 4448 35308 4768 36820
rect 10444 41972 10500 41982
rect 10444 35924 10500 41916
rect 10556 37492 10612 46172
rect 15484 46228 15540 46238
rect 11228 45332 11284 45342
rect 11228 40068 11284 45276
rect 11228 40002 11284 40012
rect 12124 43428 12180 43438
rect 10556 37426 10612 37436
rect 11788 39396 11844 39406
rect 10444 35858 10500 35868
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 2044 34804 2100 34814
rect 2044 23828 2100 34748
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 3724 33460 3780 33470
rect 2156 30996 2212 31006
rect 2156 27300 2212 30940
rect 2268 28868 2324 28878
rect 2268 28420 2324 28812
rect 2268 28354 2324 28364
rect 2156 27234 2212 27244
rect 3724 27300 3780 33404
rect 3724 27234 3780 27244
rect 4448 32172 4768 33684
rect 10332 35252 10388 35262
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 2044 23762 2100 23772
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 9100 32676 9156 32686
rect 9100 25508 9156 32620
rect 10332 32564 10388 35196
rect 10332 28420 10388 32508
rect 11676 30436 11732 30446
rect 11676 29876 11732 30380
rect 11676 29810 11732 29820
rect 10332 28354 10388 28364
rect 11788 26852 11844 39340
rect 12124 27860 12180 43372
rect 12460 41300 12516 41310
rect 12124 27794 12180 27804
rect 12236 34132 12292 34142
rect 11788 26786 11844 26796
rect 9100 25442 9156 25452
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 12236 21700 12292 34076
rect 12460 33348 12516 41244
rect 12460 32452 12516 33292
rect 12460 32386 12516 32396
rect 15036 36932 15092 36942
rect 14252 31220 14308 31230
rect 14252 28980 14308 31164
rect 15036 30548 15092 36876
rect 14252 28914 14308 28924
rect 14924 29204 14980 29214
rect 14924 28644 14980 29148
rect 14924 28578 14980 28588
rect 15036 28196 15092 30492
rect 15148 36148 15204 36158
rect 15148 28756 15204 36092
rect 15484 31780 15540 46172
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 16940 44436 16996 44446
rect 16380 44324 16436 44334
rect 15932 40740 15988 40750
rect 15484 31714 15540 31724
rect 15708 38724 15764 38734
rect 15708 29652 15764 38668
rect 15932 38668 15988 40684
rect 15932 38612 16324 38668
rect 16268 36260 16324 38612
rect 16380 37044 16436 44268
rect 16828 37828 16884 37838
rect 16380 36978 16436 36988
rect 16604 37044 16660 37054
rect 16268 30324 16324 36204
rect 16604 33572 16660 36988
rect 16604 33506 16660 33516
rect 16716 33124 16772 33134
rect 16716 31332 16772 33068
rect 16716 31266 16772 31276
rect 16268 30258 16324 30268
rect 15708 29586 15764 29596
rect 15148 28690 15204 28700
rect 15036 28130 15092 28140
rect 16828 24276 16884 37772
rect 16940 34916 16996 44380
rect 16940 34850 16996 34860
rect 18060 44324 18116 44334
rect 18060 34678 18116 44268
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19180 40628 19236 40638
rect 18172 39060 18228 39070
rect 18172 37828 18228 39004
rect 18172 37762 18228 37772
rect 18396 38612 18452 38622
rect 18060 34622 18228 34678
rect 17948 33572 18004 33582
rect 17948 29652 18004 33516
rect 18172 30884 18228 34622
rect 18396 30996 18452 38556
rect 18508 38500 18564 38510
rect 18508 37604 18564 38444
rect 18508 37538 18564 37548
rect 19180 35364 19236 40572
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19292 38612 19348 38622
rect 19292 38052 19348 38556
rect 19292 37986 19348 37996
rect 19808 37660 20128 39172
rect 19404 37604 19460 37614
rect 19404 37156 19460 37548
rect 19404 37090 19460 37100
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19180 35298 19236 35308
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19628 34916 19684 34926
rect 19628 33460 19684 34860
rect 19628 33394 19684 33404
rect 19808 34524 20128 36036
rect 20972 45444 21028 45454
rect 20412 35700 20468 35710
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 20300 34916 20356 34926
rect 19808 32956 20128 34468
rect 20188 34468 20244 34478
rect 20188 33124 20244 34412
rect 20300 33684 20356 34860
rect 20412 34580 20468 35644
rect 20412 34514 20468 34524
rect 20300 33618 20356 33628
rect 20972 33684 21028 45388
rect 25116 44996 25172 45006
rect 25116 44212 25172 44940
rect 24444 43092 24500 43102
rect 24220 42756 24276 42766
rect 20972 33618 21028 33628
rect 21084 42084 21140 42094
rect 20188 33058 20244 33068
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 18396 30930 18452 30940
rect 19516 32228 19572 32238
rect 18172 30818 18228 30828
rect 17948 29586 18004 29596
rect 18844 28868 18900 28878
rect 18844 25396 18900 28812
rect 19516 28868 19572 32172
rect 19516 28802 19572 28812
rect 19628 32004 19684 32014
rect 19628 30324 19684 31948
rect 19628 26068 19684 30268
rect 19628 26002 19684 26012
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 20412 30100 20468 30110
rect 20412 29540 20468 30044
rect 20412 29474 20468 29484
rect 20860 29876 20916 29886
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 18844 25330 18900 25340
rect 16828 24210 16884 24220
rect 19068 25284 19124 25294
rect 19068 23044 19124 25228
rect 19068 22978 19124 22988
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 20860 28980 20916 29820
rect 20860 24836 20916 28924
rect 21084 26908 21140 42028
rect 21420 41188 21476 41198
rect 21420 33908 21476 41132
rect 23100 40404 23156 40414
rect 21420 33842 21476 33852
rect 21532 39172 21588 39182
rect 20972 26852 21140 26908
rect 21420 32116 21476 32126
rect 20972 25508 21028 26852
rect 21420 26516 21476 32060
rect 21420 25732 21476 26460
rect 21420 25666 21476 25676
rect 20972 25442 21028 25452
rect 20860 24770 20916 24780
rect 21532 24052 21588 39116
rect 22876 37044 22932 37054
rect 22876 34692 22932 36988
rect 22876 34626 22932 34636
rect 23100 32452 23156 40348
rect 24220 36596 24276 42700
rect 24220 36530 24276 36540
rect 24444 36596 24500 43036
rect 25116 37380 25172 44156
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 26124 40740 26180 40750
rect 26124 39844 26180 40684
rect 26124 39778 26180 39788
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 31612 39060 31668 39070
rect 25116 37314 25172 37324
rect 28140 38612 28196 38622
rect 24444 36530 24500 36540
rect 27804 35700 27860 35710
rect 23100 32386 23156 32396
rect 23772 34804 23828 34814
rect 23772 28084 23828 34748
rect 27132 34692 27188 34702
rect 27132 31332 27188 34636
rect 27132 31266 27188 31276
rect 23772 28018 23828 28028
rect 21532 23986 21588 23996
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 12236 21634 12292 21644
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 20412 20128 21924
rect 27804 21700 27860 35644
rect 28028 35364 28084 35374
rect 28028 28532 28084 35308
rect 28028 28466 28084 28476
rect 28140 21812 28196 38556
rect 31612 38388 31668 39004
rect 31612 38322 31668 38332
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 30044 34804 30100 34814
rect 30044 27524 30100 34748
rect 30044 27458 30100 27468
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 28140 21746 28196 21756
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 27804 21634 27860 21644
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0563_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0564_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36064 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0565_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 42112 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0566_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38080 0 1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0567_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 38640 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0568_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 40096 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0569_
timestamp 1698175906
transform 1 0 32480 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0570_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39200 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0571_
timestamp 1698175906
transform -1 0 37408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0572_
timestamp 1698175906
transform -1 0 40432 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0573_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0574_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7280 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0575_
timestamp 1698175906
transform -1 0 6832 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0576_
timestamp 1698175906
transform 1 0 7392 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0577_
timestamp 1698175906
transform -1 0 9184 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0578_
timestamp 1698175906
transform 1 0 3360 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0579_
timestamp 1698175906
transform 1 0 8064 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0580_
timestamp 1698175906
transform 1 0 2016 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0581_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4368 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0582_
timestamp 1698175906
transform 1 0 9520 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0583_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0584_
timestamp 1698175906
transform -1 0 15456 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0585_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28448 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0586_
timestamp 1698175906
transform 1 0 39088 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0587_
timestamp 1698175906
transform -1 0 37744 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0588_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0589_
timestamp 1698175906
transform -1 0 39760 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _0590_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32704 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0591_
timestamp 1698175906
transform 1 0 41328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0592_
timestamp 1698175906
transform -1 0 35056 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0593_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 34384 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0594_
timestamp 1698175906
transform -1 0 31136 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0595_
timestamp 1698175906
transform 1 0 2800 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0596_
timestamp 1698175906
transform 1 0 3360 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0597_
timestamp 1698175906
transform 1 0 3808 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0598_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7392 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0599_
timestamp 1698175906
transform 1 0 7952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0600_
timestamp 1698175906
transform -1 0 10192 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0601_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6944 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0602_
timestamp 1698175906
transform -1 0 7952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0603_
timestamp 1698175906
transform -1 0 12320 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0604_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0605_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0606_
timestamp 1698175906
transform 1 0 14112 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0607_
timestamp 1698175906
transform -1 0 6944 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0608_
timestamp 1698175906
transform -1 0 7392 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0609_
timestamp 1698175906
transform -1 0 7056 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0610_
timestamp 1698175906
transform 1 0 3808 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0611_
timestamp 1698175906
transform -1 0 9184 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0612_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13552 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0613_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3248 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0614_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6384 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0615_
timestamp 1698175906
transform -1 0 6384 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0616_
timestamp 1698175906
transform 1 0 13776 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0617_
timestamp 1698175906
transform -1 0 39088 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0618_
timestamp 1698175906
transform 1 0 37184 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0619_
timestamp 1698175906
transform -1 0 12656 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0620_
timestamp 1698175906
transform -1 0 12656 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0621_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 39200 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0622_
timestamp 1698175906
transform -1 0 36400 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0623_
timestamp 1698175906
transform -1 0 35168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0624_
timestamp 1698175906
transform 1 0 32704 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0625_
timestamp 1698175906
transform -1 0 32368 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0626_
timestamp 1698175906
transform 1 0 2912 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0627_
timestamp 1698175906
transform -1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _0628_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11648 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0629_
timestamp 1698175906
transform -1 0 7840 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0630_
timestamp 1698175906
transform -1 0 8064 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0631_
timestamp 1698175906
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0632_
timestamp 1698175906
transform -1 0 9856 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0633_
timestamp 1698175906
transform -1 0 33712 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0634_
timestamp 1698175906
transform -1 0 32480 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0635_
timestamp 1698175906
transform -1 0 32704 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0636_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32256 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0637_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19264 0 1 39200
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0638_
timestamp 1698175906
transform 1 0 15008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0639_
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0640_
timestamp 1698175906
transform 1 0 36960 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0641_
timestamp 1698175906
transform -1 0 38864 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0642_
timestamp 1698175906
transform 1 0 34048 0 -1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0643_
timestamp 1698175906
transform -1 0 31024 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0644_
timestamp 1698175906
transform 1 0 28112 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0645_
timestamp 1698175906
transform 1 0 21168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0646_
timestamp 1698175906
transform 1 0 37408 0 1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0647_
timestamp 1698175906
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0648_
timestamp 1698175906
transform -1 0 40992 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0649_
timestamp 1698175906
transform -1 0 31360 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0650_
timestamp 1698175906
transform 1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0651_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5712 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0652_
timestamp 1698175906
transform -1 0 8064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0653_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23072 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0654_
timestamp 1698175906
transform -1 0 36624 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0655_
timestamp 1698175906
transform -1 0 31136 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0656_
timestamp 1698175906
transform 1 0 34496 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0657_
timestamp 1698175906
transform 1 0 27664 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0658_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11648 0 -1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0659_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28224 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0660_
timestamp 1698175906
transform -1 0 10976 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0661_
timestamp 1698175906
transform 1 0 22064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0662_
timestamp 1698175906
transform -1 0 7840 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0663_
timestamp 1698175906
transform 1 0 14112 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0664_
timestamp 1698175906
transform -1 0 30688 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0665_
timestamp 1698175906
transform 1 0 28672 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0666_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0667_
timestamp 1698175906
transform 1 0 10192 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0668_
timestamp 1698175906
transform 1 0 14224 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0669_
timestamp 1698175906
transform 1 0 22288 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0670_
timestamp 1698175906
transform 1 0 6384 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0671_
timestamp 1698175906
transform 1 0 8624 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0672_
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0673_
timestamp 1698175906
transform -1 0 36624 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0674_
timestamp 1698175906
transform -1 0 25984 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0675_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28112 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0676_
timestamp 1698175906
transform -1 0 31584 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0677_
timestamp 1698175906
transform 1 0 11648 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0678_
timestamp 1698175906
transform 1 0 7504 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0679_
timestamp 1698175906
transform 1 0 20272 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0680_
timestamp 1698175906
transform -1 0 26320 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0681_
timestamp 1698175906
transform -1 0 24528 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0682_
timestamp 1698175906
transform 1 0 24752 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0683_
timestamp 1698175906
transform 1 0 25200 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0684_
timestamp 1698175906
transform -1 0 10976 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0685_
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0686_
timestamp 1698175906
transform 1 0 11984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0687_
timestamp 1698175906
transform 1 0 6720 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0688_
timestamp 1698175906
transform 1 0 7952 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0689_
timestamp 1698175906
transform 1 0 9520 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0690_
timestamp 1698175906
transform 1 0 9632 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0691_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13104 0 -1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0692_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0693_
timestamp 1698175906
transform 1 0 13328 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0694_
timestamp 1698175906
transform -1 0 16688 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0695_
timestamp 1698175906
transform -1 0 9184 0 -1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0696_
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0697_
timestamp 1698175906
transform -1 0 37072 0 -1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0698_
timestamp 1698175906
transform -1 0 24080 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0699_
timestamp 1698175906
transform -1 0 8736 0 1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0700_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16912 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0701_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14560 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0702_
timestamp 1698175906
transform -1 0 13888 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0703_
timestamp 1698175906
transform -1 0 34384 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0704_
timestamp 1698175906
transform -1 0 21952 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0705_
timestamp 1698175906
transform -1 0 4480 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _0706_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6384 0 1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0707_
timestamp 1698175906
transform -1 0 10752 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0708_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 38640 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0709_
timestamp 1698175906
transform -1 0 4032 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0710_
timestamp 1698175906
transform 1 0 5376 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0711_
timestamp 1698175906
transform -1 0 4144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0712_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6048 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0713_
timestamp 1698175906
transform -1 0 9184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0714_
timestamp 1698175906
transform -1 0 32256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0715_
timestamp 1698175906
transform 1 0 6048 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0716_
timestamp 1698175906
transform -1 0 7952 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0717_
timestamp 1698175906
transform -1 0 12096 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0718_
timestamp 1698175906
transform -1 0 12320 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0719_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0720_
timestamp 1698175906
transform -1 0 20272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0721_
timestamp 1698175906
transform -1 0 18368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0722_
timestamp 1698175906
transform 1 0 32144 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0723_
timestamp 1698175906
transform -1 0 23968 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0724_
timestamp 1698175906
transform 1 0 22848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0725_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17696 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0726_
timestamp 1698175906
transform 1 0 17360 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0727_
timestamp 1698175906
transform -1 0 24976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0728_
timestamp 1698175906
transform -1 0 24080 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0729_
timestamp 1698175906
transform 1 0 15568 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0730_
timestamp 1698175906
transform 1 0 13664 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0731_
timestamp 1698175906
transform -1 0 30128 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0732_
timestamp 1698175906
transform -1 0 6384 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0733_
timestamp 1698175906
transform -1 0 16352 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0734_
timestamp 1698175906
transform 1 0 15120 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0735_
timestamp 1698175906
transform -1 0 3248 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0736_
timestamp 1698175906
transform -1 0 3584 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0737_
timestamp 1698175906
transform 1 0 3472 0 -1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0738_
timestamp 1698175906
transform -1 0 3248 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0739_
timestamp 1698175906
transform 1 0 33712 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0740_
timestamp 1698175906
transform -1 0 35840 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0741_
timestamp 1698175906
transform 1 0 11760 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0742_
timestamp 1698175906
transform 1 0 33600 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _0743_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27888 0 -1 40768
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0744_
timestamp 1698175906
transform 1 0 2128 0 -1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0745_
timestamp 1698175906
transform -1 0 12320 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0746_
timestamp 1698175906
transform 1 0 5712 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0747_
timestamp 1698175906
transform -1 0 5264 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0748_
timestamp 1698175906
transform 1 0 3248 0 1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0749_
timestamp 1698175906
transform -1 0 2912 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0750_
timestamp 1698175906
transform 1 0 2352 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0751_
timestamp 1698175906
transform 1 0 4144 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0752_
timestamp 1698175906
transform -1 0 10640 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0753_
timestamp 1698175906
transform -1 0 9184 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0754_
timestamp 1698175906
transform 1 0 13328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0755_
timestamp 1698175906
transform -1 0 12992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0756_
timestamp 1698175906
transform 1 0 9968 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0757_
timestamp 1698175906
transform -1 0 14896 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0758_
timestamp 1698175906
transform -1 0 9296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0759_
timestamp 1698175906
transform -1 0 14224 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0760_
timestamp 1698175906
transform -1 0 12992 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0761_
timestamp 1698175906
transform -1 0 9408 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0762_
timestamp 1698175906
transform 1 0 15456 0 1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0763_
timestamp 1698175906
transform -1 0 19152 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0764_
timestamp 1698175906
transform -1 0 19376 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0765_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 -1 25088
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0766_
timestamp 1698175906
transform 1 0 21168 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0767_
timestamp 1698175906
transform 1 0 13776 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0768_
timestamp 1698175906
transform -1 0 15792 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0769_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22848 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0770_
timestamp 1698175906
transform 1 0 13552 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0771_
timestamp 1698175906
transform 1 0 19264 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0772_
timestamp 1698175906
transform -1 0 21280 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0773_
timestamp 1698175906
transform 1 0 7952 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0774_
timestamp 1698175906
transform 1 0 22064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0775_
timestamp 1698175906
transform 1 0 20272 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0776_
timestamp 1698175906
transform 1 0 5600 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0777_
timestamp 1698175906
transform 1 0 21504 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0778_
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0779_
timestamp 1698175906
transform -1 0 26880 0 1 25088
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0780_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8288 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0781_
timestamp 1698175906
transform -1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0782_
timestamp 1698175906
transform 1 0 30240 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0783_
timestamp 1698175906
transform -1 0 27328 0 1 36064
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0784_
timestamp 1698175906
transform -1 0 24864 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0785_
timestamp 1698175906
transform 1 0 7504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0786_
timestamp 1698175906
transform 1 0 20048 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0787_
timestamp 1698175906
transform -1 0 31136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _0788_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 -1 34496
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0789_
timestamp 1698175906
transform -1 0 20272 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0790_
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0791_
timestamp 1698175906
transform -1 0 29904 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0792_
timestamp 1698175906
transform 1 0 18256 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0793_
timestamp 1698175906
transform 1 0 19600 0 -1 37632
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0794_
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0795_
timestamp 1698175906
transform 1 0 23968 0 1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0796_
timestamp 1698175906
transform 1 0 7840 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0797_
timestamp 1698175906
transform 1 0 11648 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0798_
timestamp 1698175906
transform -1 0 27888 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0799_
timestamp 1698175906
transform -1 0 25648 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0800_
timestamp 1698175906
transform -1 0 28000 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0801_
timestamp 1698175906
transform -1 0 26656 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0802_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8064 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0803_
timestamp 1698175906
transform -1 0 9184 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0804_
timestamp 1698175906
transform 1 0 9296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0805_
timestamp 1698175906
transform -1 0 13104 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0806_
timestamp 1698175906
transform 1 0 9520 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0807_
timestamp 1698175906
transform 1 0 9184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0808_
timestamp 1698175906
transform -1 0 11648 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0809_
timestamp 1698175906
transform 1 0 11648 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0810_
timestamp 1698175906
transform 1 0 10192 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0811_
timestamp 1698175906
transform 1 0 23296 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0812_
timestamp 1698175906
transform -1 0 27216 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0813_
timestamp 1698175906
transform 1 0 25200 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0814_
timestamp 1698175906
transform 1 0 26320 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0815_
timestamp 1698175906
transform 1 0 26096 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0816_
timestamp 1698175906
transform 1 0 24976 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0817_
timestamp 1698175906
transform 1 0 15792 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0818_
timestamp 1698175906
transform 1 0 13440 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0819_
timestamp 1698175906
transform -1 0 26768 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0820_
timestamp 1698175906
transform -1 0 18928 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0821_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15792 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0822_
timestamp 1698175906
transform -1 0 20160 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0823_
timestamp 1698175906
transform -1 0 17696 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0824_
timestamp 1698175906
transform 1 0 17024 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0825_
timestamp 1698175906
transform -1 0 23184 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0826_
timestamp 1698175906
transform -1 0 18704 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0827_
timestamp 1698175906
transform -1 0 16128 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0828_
timestamp 1698175906
transform 1 0 17248 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0829_
timestamp 1698175906
transform -1 0 4144 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0830_
timestamp 1698175906
transform 1 0 2128 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0831_
timestamp 1698175906
transform 1 0 3584 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0832_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _0833_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0834_
timestamp 1698175906
transform 1 0 12992 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0835_
timestamp 1698175906
transform 1 0 14448 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0836_
timestamp 1698175906
transform 1 0 16016 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0837_
timestamp 1698175906
transform 1 0 17472 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0838_
timestamp 1698175906
transform 1 0 16464 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0839_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0840_
timestamp 1698175906
transform 1 0 16016 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0841_
timestamp 1698175906
transform -1 0 32480 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0842_
timestamp 1698175906
transform -1 0 30240 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0843_
timestamp 1698175906
transform 1 0 28224 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0844_
timestamp 1698175906
transform -1 0 30800 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0845_
timestamp 1698175906
transform 1 0 10416 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0846_
timestamp 1698175906
transform 1 0 12768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0847_
timestamp 1698175906
transform 1 0 21504 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0848_
timestamp 1698175906
transform -1 0 24864 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0849_
timestamp 1698175906
transform 1 0 23520 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0850_
timestamp 1698175906
transform -1 0 12656 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0851_
timestamp 1698175906
transform -1 0 28560 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0852_
timestamp 1698175906
transform 1 0 11536 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0853_
timestamp 1698175906
transform 1 0 12544 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0854_
timestamp 1698175906
transform -1 0 14336 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0855_
timestamp 1698175906
transform -1 0 26432 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0856_
timestamp 1698175906
transform 1 0 25984 0 -1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0857_
timestamp 1698175906
transform 1 0 26768 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0858_
timestamp 1698175906
transform 1 0 24416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0859_
timestamp 1698175906
transform -1 0 23520 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0860_
timestamp 1698175906
transform -1 0 26544 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0861_
timestamp 1698175906
transform 1 0 27440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0862_
timestamp 1698175906
transform -1 0 28448 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0863_
timestamp 1698175906
transform -1 0 29568 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0864_
timestamp 1698175906
transform -1 0 28784 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0865_
timestamp 1698175906
transform -1 0 3808 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0866_
timestamp 1698175906
transform 1 0 1792 0 -1 32928
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0867_
timestamp 1698175906
transform 1 0 5264 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0868_
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0869_
timestamp 1698175906
transform -1 0 19264 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0870_
timestamp 1698175906
transform 1 0 12768 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0871_
timestamp 1698175906
transform 1 0 2352 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0872_
timestamp 1698175906
transform 1 0 15904 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0873_
timestamp 1698175906
transform -1 0 17808 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0874_
timestamp 1698175906
transform 1 0 17024 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0875_
timestamp 1698175906
transform 1 0 17360 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0876_
timestamp 1698175906
transform 1 0 25760 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0877_
timestamp 1698175906
transform -1 0 19040 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0878_
timestamp 1698175906
transform -1 0 21840 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0879_
timestamp 1698175906
transform -1 0 22736 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0880_
timestamp 1698175906
transform 1 0 18256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0881_
timestamp 1698175906
transform -1 0 26208 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0882_
timestamp 1698175906
transform -1 0 10304 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0883_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0884_
timestamp 1698175906
transform 1 0 17584 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0885_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18144 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0886_
timestamp 1698175906
transform 1 0 9632 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0887_
timestamp 1698175906
transform 1 0 17696 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0888_
timestamp 1698175906
transform -1 0 20160 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0889_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0890_
timestamp 1698175906
transform 1 0 18032 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0891_
timestamp 1698175906
transform -1 0 18480 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0892_
timestamp 1698175906
transform 1 0 18256 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0893_
timestamp 1698175906
transform 1 0 18368 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0894_
timestamp 1698175906
transform -1 0 24640 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0895_
timestamp 1698175906
transform -1 0 30016 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0896_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26320 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0897_
timestamp 1698175906
transform -1 0 28672 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0898_
timestamp 1698175906
transform -1 0 19264 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0899_
timestamp 1698175906
transform -1 0 28112 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0900_
timestamp 1698175906
transform 1 0 27104 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0901_
timestamp 1698175906
transform -1 0 28000 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0902_
timestamp 1698175906
transform -1 0 6272 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0903_
timestamp 1698175906
transform 1 0 8176 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0904_
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0905_
timestamp 1698175906
transform 1 0 7840 0 1 31360
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0906_
timestamp 1698175906
transform -1 0 14112 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0907_
timestamp 1698175906
transform 1 0 14560 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0908_
timestamp 1698175906
transform 1 0 13776 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0909_
timestamp 1698175906
transform 1 0 14224 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0910_
timestamp 1698175906
transform 1 0 23072 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0911_
timestamp 1698175906
transform 1 0 13776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0912_
timestamp 1698175906
transform 1 0 21392 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0913_
timestamp 1698175906
transform 1 0 22736 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0914_
timestamp 1698175906
transform 1 0 23744 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0915_
timestamp 1698175906
transform 1 0 24640 0 1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0916_
timestamp 1698175906
transform 1 0 24864 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0917_
timestamp 1698175906
transform 1 0 27440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0918_
timestamp 1698175906
transform 1 0 28112 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0919_
timestamp 1698175906
transform 1 0 24416 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0920_
timestamp 1698175906
transform 1 0 26432 0 -1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0921_
timestamp 1698175906
transform -1 0 26096 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0922_
timestamp 1698175906
transform -1 0 26096 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0923_
timestamp 1698175906
transform 1 0 18368 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0924_
timestamp 1698175906
transform -1 0 26880 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0925_
timestamp 1698175906
transform -1 0 26768 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0926_
timestamp 1698175906
transform -1 0 25984 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0927_
timestamp 1698175906
transform 1 0 23296 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0928_
timestamp 1698175906
transform -1 0 10864 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0929_
timestamp 1698175906
transform -1 0 9184 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0930_
timestamp 1698175906
transform -1 0 11424 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0931_
timestamp 1698175906
transform -1 0 11200 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0932_
timestamp 1698175906
transform -1 0 8960 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0933_
timestamp 1698175906
transform 1 0 1904 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0934_
timestamp 1698175906
transform 1 0 3696 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0935_
timestamp 1698175906
transform 1 0 2240 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0936_
timestamp 1698175906
transform 1 0 2912 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0937_
timestamp 1698175906
transform -1 0 14560 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0938_
timestamp 1698175906
transform -1 0 21952 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0939_
timestamp 1698175906
transform 1 0 8960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0940_
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0941_
timestamp 1698175906
transform -1 0 5600 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0942_
timestamp 1698175906
transform 1 0 5600 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0943_
timestamp 1698175906
transform 1 0 6272 0 1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0944_
timestamp 1698175906
transform 1 0 17248 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0945_
timestamp 1698175906
transform -1 0 21840 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0946_
timestamp 1698175906
transform 1 0 22512 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0947_
timestamp 1698175906
transform 1 0 17360 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0948_
timestamp 1698175906
transform 1 0 19488 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0949_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22736 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0950_
timestamp 1698175906
transform 1 0 25200 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0951_
timestamp 1698175906
transform 1 0 29008 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0952_
timestamp 1698175906
transform -1 0 38976 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0953_
timestamp 1698175906
transform 1 0 29008 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0954_
timestamp 1698175906
transform -1 0 22624 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0955_
timestamp 1698175906
transform 1 0 20160 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0956_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0957_
timestamp 1698175906
transform 1 0 18592 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0958_
timestamp 1698175906
transform -1 0 19712 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0959_
timestamp 1698175906
transform 1 0 15232 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0960_
timestamp 1698175906
transform 1 0 15680 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0961_
timestamp 1698175906
transform -1 0 4368 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0962_
timestamp 1698175906
transform 1 0 2352 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0963_
timestamp 1698175906
transform 1 0 2128 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0964_
timestamp 1698175906
transform 1 0 3136 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0965_
timestamp 1698175906
transform 1 0 17472 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0966_
timestamp 1698175906
transform 1 0 22624 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0967_
timestamp 1698175906
transform -1 0 28560 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0968_
timestamp 1698175906
transform -1 0 27104 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0969_
timestamp 1698175906
transform 1 0 25984 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0970_
timestamp 1698175906
transform -1 0 31920 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0971_
timestamp 1698175906
transform 1 0 29008 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0972_
timestamp 1698175906
transform -1 0 40320 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0973_
timestamp 1698175906
transform 1 0 28112 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0974_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26544 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0975_
timestamp 1698175906
transform -1 0 20496 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0976_
timestamp 1698175906
transform -1 0 20944 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0977_
timestamp 1698175906
transform 1 0 19488 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0978_
timestamp 1698175906
transform 1 0 20832 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0979_
timestamp 1698175906
transform -1 0 11536 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _0980_
timestamp 1698175906
transform 1 0 7392 0 1 29792
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _0981_
timestamp 1698175906
transform 1 0 1792 0 1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0982_
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0983_
timestamp 1698175906
transform 1 0 26432 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0984_
timestamp 1698175906
transform 1 0 19824 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0985_
timestamp 1698175906
transform -1 0 15568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0986_
timestamp 1698175906
transform 1 0 16464 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0987_
timestamp 1698175906
transform 1 0 15344 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0988_
timestamp 1698175906
transform -1 0 21728 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0989_
timestamp 1698175906
transform -1 0 18480 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0990_
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0991_
timestamp 1698175906
transform 1 0 15008 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0992_
timestamp 1698175906
transform 1 0 16240 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0993_
timestamp 1698175906
transform 1 0 22624 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0994_
timestamp 1698175906
transform 1 0 23184 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0995_
timestamp 1698175906
transform 1 0 23184 0 1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0996_
timestamp 1698175906
transform 1 0 31024 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0997_
timestamp 1698175906
transform -1 0 38976 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _0998_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 31024 0 1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0999_
timestamp 1698175906
transform 1 0 30576 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1000_
timestamp 1698175906
transform 1 0 20384 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1001_
timestamp 1698175906
transform 1 0 18928 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1002_
timestamp 1698175906
transform 1 0 19936 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1003_
timestamp 1698175906
transform -1 0 20608 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1004_
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1005_
timestamp 1698175906
transform 1 0 21168 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1006_
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1007_
timestamp 1698175906
transform 1 0 2128 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1008_
timestamp 1698175906
transform 1 0 3136 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1009_
timestamp 1698175906
transform -1 0 9184 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1010_
timestamp 1698175906
transform 1 0 3808 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1011_
timestamp 1698175906
transform 1 0 19040 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1012_
timestamp 1698175906
transform 1 0 20160 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1013_
timestamp 1698175906
transform 1 0 20608 0 -1 47040
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1014_
timestamp 1698175906
transform 1 0 21728 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1015_
timestamp 1698175906
transform 1 0 30800 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1016_
timestamp 1698175906
transform -1 0 37632 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1017_
timestamp 1698175906
transform 1 0 27664 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1018_
timestamp 1698175906
transform -1 0 30800 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1019_
timestamp 1698175906
transform -1 0 19488 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1020_
timestamp 1698175906
transform -1 0 20720 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1021_
timestamp 1698175906
transform -1 0 20272 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1022_
timestamp 1698175906
transform 1 0 12432 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1023_
timestamp 1698175906
transform -1 0 14448 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1024_
timestamp 1698175906
transform 1 0 14560 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1025_
timestamp 1698175906
transform 1 0 15904 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1026_
timestamp 1698175906
transform 1 0 14672 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1027_
timestamp 1698175906
transform 1 0 14784 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1028_
timestamp 1698175906
transform 1 0 2128 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1029_
timestamp 1698175906
transform -1 0 3136 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1030_
timestamp 1698175906
transform 1 0 2576 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1031_
timestamp 1698175906
transform 1 0 18368 0 -1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1032_
timestamp 1698175906
transform 1 0 30464 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1033_
timestamp 1698175906
transform -1 0 23184 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1034_
timestamp 1698175906
transform -1 0 10416 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1035_
timestamp 1698175906
transform 1 0 11648 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1036_
timestamp 1698175906
transform 1 0 12992 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1037_
timestamp 1698175906
transform -1 0 12544 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1038_
timestamp 1698175906
transform 1 0 12656 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1039_
timestamp 1698175906
transform 1 0 11760 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1040_
timestamp 1698175906
transform 1 0 10528 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1041_
timestamp 1698175906
transform -1 0 25648 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1042_
timestamp 1698175906
transform 1 0 11088 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1043_
timestamp 1698175906
transform 1 0 9856 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1044_
timestamp 1698175906
transform -1 0 27888 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698175906
transform 1 0 10976 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1046_
timestamp 1698175906
transform 1 0 10416 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1047_
timestamp 1698175906
transform -1 0 29792 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1048_
timestamp 1698175906
transform 1 0 31584 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1049_
timestamp 1698175906
transform 1 0 12320 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1050_
timestamp 1698175906
transform 1 0 10976 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1051_
timestamp 1698175906
transform -1 0 32928 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1052_
timestamp 1698175906
transform 1 0 32928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1053_
timestamp 1698175906
transform -1 0 35504 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1054_
timestamp 1698175906
transform 1 0 35840 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1055_
timestamp 1698175906
transform 1 0 34944 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1056_
timestamp 1698175906
transform -1 0 35168 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1057_
timestamp 1698175906
transform 1 0 34160 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1058_
timestamp 1698175906
transform 1 0 34720 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1059_
timestamp 1698175906
transform 1 0 36848 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1060_
timestamp 1698175906
transform 1 0 34160 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1061_
timestamp 1698175906
transform 1 0 34832 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1062_
timestamp 1698175906
transform -1 0 39312 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1063_
timestamp 1698175906
transform 1 0 33488 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1064_
timestamp 1698175906
transform -1 0 35168 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1065_
timestamp 1698175906
transform 1 0 14784 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1066_
timestamp 1698175906
transform 1 0 21952 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1067_
timestamp 1698175906
transform -1 0 25984 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1068_
timestamp 1698175906
transform 1 0 12320 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1069_
timestamp 1698175906
transform -1 0 27216 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1070_
timestamp 1698175906
transform 1 0 24416 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1071_
timestamp 1698175906
transform 1 0 22288 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1072_
timestamp 1698175906
transform 1 0 26096 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1073_
timestamp 1698175906
transform 1 0 24416 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1074_
timestamp 1698175906
transform 1 0 23408 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1075_
timestamp 1698175906
transform 1 0 22176 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1076_
timestamp 1698175906
transform -1 0 26320 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1077_
timestamp 1698175906
transform 1 0 26208 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1078_
timestamp 1698175906
transform 1 0 38640 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1079_
timestamp 1698175906
transform 1 0 38976 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1080_
timestamp 1698175906
transform 1 0 38304 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1081_
timestamp 1698175906
transform -1 0 39872 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1082_
timestamp 1698175906
transform -1 0 41664 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1083_
timestamp 1698175906
transform 1 0 40992 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1084_
timestamp 1698175906
transform 1 0 40320 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1085_
timestamp 1698175906
transform -1 0 39872 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1086_
timestamp 1698175906
transform 1 0 38864 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1087_
timestamp 1698175906
transform -1 0 41440 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1088_
timestamp 1698175906
transform -1 0 42112 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1089_
timestamp 1698175906
transform 1 0 29008 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1090_
timestamp 1698175906
transform 1 0 32816 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1091_
timestamp 1698175906
transform -1 0 38640 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1092_
timestamp 1698175906
transform -1 0 32256 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1093_
timestamp 1698175906
transform 1 0 29680 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1094_
timestamp 1698175906
transform -1 0 32368 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1095_
timestamp 1698175906
transform 1 0 29792 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1096_
timestamp 1698175906
transform -1 0 36624 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1097_
timestamp 1698175906
transform 1 0 33040 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1098_
timestamp 1698175906
transform -1 0 38528 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1099_
timestamp 1698175906
transform 1 0 36848 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1100_
timestamp 1698175906
transform 1 0 32928 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1101_
timestamp 1698175906
transform 1 0 39088 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1102_
timestamp 1698175906
transform 1 0 38416 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1103_
timestamp 1698175906
transform -1 0 40544 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1104_
timestamp 1698175906
transform -1 0 39872 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1105_
timestamp 1698175906
transform -1 0 42560 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1106_
timestamp 1698175906
transform 1 0 40768 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1107_
timestamp 1698175906
transform -1 0 42672 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1108_
timestamp 1698175906
transform 1 0 40880 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1109_
timestamp 1698175906
transform 1 0 40768 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1110_
timestamp 1698175906
transform 1 0 40768 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1111_
timestamp 1698175906
transform 1 0 15008 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1112_
timestamp 1698175906
transform -1 0 17024 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1113_
timestamp 1698175906
transform 1 0 17248 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1114_
timestamp 1698175906
transform 1 0 16128 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1115_
timestamp 1698175906
transform 1 0 15568 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1116_
timestamp 1698175906
transform 1 0 14448 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1117_
timestamp 1698175906
transform 1 0 15344 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1118_
timestamp 1698175906
transform 1 0 14448 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1119_
timestamp 1698175906
transform 1 0 18144 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1120_
timestamp 1698175906
transform 1 0 17248 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1121_
timestamp 1698175906
transform 1 0 18032 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1122_
timestamp 1698175906
transform 1 0 17920 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1123_
timestamp 1698175906
transform 1 0 30352 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1124_
timestamp 1698175906
transform 1 0 30128 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1125_
timestamp 1698175906
transform -1 0 33936 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1126_
timestamp 1698175906
transform 1 0 32592 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1127_
timestamp 1698175906
transform -1 0 33824 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1128_
timestamp 1698175906
transform 1 0 34048 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1129_
timestamp 1698175906
transform -1 0 35840 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1130_
timestamp 1698175906
transform 1 0 34160 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1131_
timestamp 1698175906
transform -1 0 35392 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1132_
timestamp 1698175906
transform 1 0 32704 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1133_
timestamp 1698175906
transform 1 0 31024 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1134_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4816 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1135_
timestamp 1698175906
transform -1 0 4816 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1136_
timestamp 1698175906
transform -1 0 8960 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1137_
timestamp 1698175906
transform 1 0 4144 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1138_
timestamp 1698175906
transform 1 0 36848 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1139_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 35056 0 -1 37632
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1140_
timestamp 1698175906
transform 1 0 37296 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1141_
timestamp 1698175906
transform 1 0 33712 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1142_
timestamp 1698175906
transform 1 0 21168 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1143_
timestamp 1698175906
transform 1 0 25088 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1144_
timestamp 1698175906
transform 1 0 20832 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1145_
timestamp 1698175906
transform 1 0 25200 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1146_
timestamp 1698175906
transform -1 0 43120 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1147_
timestamp 1698175906
transform 1 0 40768 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1148_
timestamp 1698175906
transform -1 0 40320 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1149_
timestamp 1698175906
transform 1 0 41440 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1150_
timestamp 1698175906
transform 1 0 29008 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1151_
timestamp 1698175906
transform 1 0 29232 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1152_
timestamp 1698175906
transform 1 0 33376 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1153_
timestamp 1698175906
transform 1 0 33152 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1154_
timestamp 1698175906
transform 1 0 37072 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1155_
timestamp 1698175906
transform 1 0 41888 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1156_
timestamp 1698175906
transform 1 0 41104 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1157_
timestamp 1698175906
transform 1 0 40096 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1158_
timestamp 1698175906
transform 1 0 13328 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1159_
timestamp 1698175906
transform 1 0 12992 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1160_
timestamp 1698175906
transform 1 0 17472 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1161_
timestamp 1698175906
transform -1 0 20944 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1162_
timestamp 1698175906
transform -1 0 32704 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1163_
timestamp 1698175906
transform -1 0 37520 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1164_
timestamp 1698175906
transform -1 0 37632 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1165_
timestamp 1698175906
transform -1 0 32368 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__A1 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__A2
timestamp 1698175906
transform 1 0 15680 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0585__I
timestamp 1698175906
transform 1 0 24752 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0612__A3
timestamp 1698175906
transform 1 0 15120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0619__I
timestamp 1698175906
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__A3
timestamp 1698175906
transform -1 0 29680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__B1
timestamp 1698175906
transform -1 0 29680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0637__A1
timestamp 1698175906
transform -1 0 19712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0637__B1
timestamp 1698175906
transform -1 0 14784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0637__B2
timestamp 1698175906
transform 1 0 14112 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0644__A1
timestamp 1698175906
transform 1 0 27440 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0644__A2
timestamp 1698175906
transform -1 0 28112 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0647__I
timestamp 1698175906
transform 1 0 26208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__A1
timestamp 1698175906
transform -1 0 23072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__B1
timestamp 1698175906
transform 1 0 25088 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__B2
timestamp 1698175906
transform 1 0 22624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0657__I
timestamp 1698175906
transform 1 0 29232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0659__A1
timestamp 1698175906
transform -1 0 27328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0659__A2
timestamp 1698175906
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0659__B
timestamp 1698175906
transform 1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0665__A2
timestamp 1698175906
transform 1 0 28448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0668__I
timestamp 1698175906
transform 1 0 14000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0669__A1
timestamp 1698175906
transform -1 0 23520 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0674__I
timestamp 1698175906
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0675__A1
timestamp 1698175906
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0675__A2
timestamp 1698175906
transform -1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0677__I
timestamp 1698175906
transform 1 0 12544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0679__A1
timestamp 1698175906
transform 1 0 20048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0680__I
timestamp 1698175906
transform 1 0 26544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0681__A1
timestamp 1698175906
transform 1 0 23744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0683__A2
timestamp 1698175906
transform 1 0 27552 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0686__I
timestamp 1698175906
transform 1 0 13552 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0692__B2
timestamp 1698175906
transform 1 0 14448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0693__A1
timestamp 1698175906
transform 1 0 16240 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0693__A2
timestamp 1698175906
transform 1 0 16464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0699__B
timestamp 1698175906
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0700__A3
timestamp 1698175906
transform -1 0 15456 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0701__A1
timestamp 1698175906
transform 1 0 15232 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0701__A2
timestamp 1698175906
transform -1 0 15008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0704__I
timestamp 1698175906
transform 1 0 22176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0706__A2
timestamp 1698175906
transform -1 0 6384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0709__I
timestamp 1698175906
transform 1 0 4256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0716__I
timestamp 1698175906
transform 1 0 6832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0718__A2
timestamp 1698175906
transform -1 0 11760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0718__B1
timestamp 1698175906
transform -1 0 11312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0719__A1
timestamp 1698175906
transform 1 0 12544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0723__I
timestamp 1698175906
transform -1 0 24192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0726__A3
timestamp 1698175906
transform 1 0 21392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__I
timestamp 1698175906
transform -1 0 25536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0729__A2
timestamp 1698175906
transform -1 0 14784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0733__A2
timestamp 1698175906
transform -1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0733__B1
timestamp 1698175906
transform 1 0 14112 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0733__B2
timestamp 1698175906
transform 1 0 16352 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0735__A1
timestamp 1698175906
transform -1 0 3472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0737__A4
timestamp 1698175906
transform 1 0 6048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__A3
timestamp 1698175906
transform 1 0 27216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__B2
timestamp 1698175906
transform -1 0 27888 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0744__A1
timestamp 1698175906
transform 1 0 6048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0744__C
timestamp 1698175906
transform 1 0 5824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0745__A2
timestamp 1698175906
transform 1 0 12992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__A1
timestamp 1698175906
transform -1 0 4704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__A2
timestamp 1698175906
transform -1 0 4256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0748__A3
timestamp 1698175906
transform 1 0 5152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0752__I
timestamp 1698175906
transform 1 0 10640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0755__I
timestamp 1698175906
transform 1 0 13216 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0756__A2
timestamp 1698175906
transform -1 0 15568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0756__B
timestamp 1698175906
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0759__I
timestamp 1698175906
transform -1 0 13776 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0761__A3
timestamp 1698175906
transform 1 0 9632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__I
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A1
timestamp 1698175906
transform -1 0 11760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A2
timestamp 1698175906
transform -1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0768__I
timestamp 1698175906
transform -1 0 15680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0769__A1
timestamp 1698175906
transform -1 0 23072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0769__A2
timestamp 1698175906
transform -1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0771__A1
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0771__A2
timestamp 1698175906
transform 1 0 19488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0771__B
timestamp 1698175906
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__I
timestamp 1698175906
transform 1 0 23184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A1
timestamp 1698175906
transform 1 0 29792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A2
timestamp 1698175906
transform -1 0 25536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__B2
timestamp 1698175906
transform -1 0 21616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0778__I
timestamp 1698175906
transform 1 0 8176 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__A1
timestamp 1698175906
transform -1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__B2
timestamp 1698175906
transform 1 0 19936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__C1
timestamp 1698175906
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__C2
timestamp 1698175906
transform 1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0780__A3
timestamp 1698175906
transform 1 0 8512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__A1
timestamp 1698175906
transform 1 0 29120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__A2
timestamp 1698175906
transform 1 0 20160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__B1
timestamp 1698175906
transform 1 0 21392 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__B2
timestamp 1698175906
transform 1 0 29680 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__C2
timestamp 1698175906
transform 1 0 21840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__A1
timestamp 1698175906
transform 1 0 19712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__A2
timestamp 1698175906
transform -1 0 22064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__B
timestamp 1698175906
transform -1 0 19488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__B1
timestamp 1698175906
transform 1 0 18032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__B2
timestamp 1698175906
transform 1 0 19488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__C1
timestamp 1698175906
transform 1 0 20272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__C2
timestamp 1698175906
transform 1 0 19488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__A1
timestamp 1698175906
transform 1 0 19376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__A2
timestamp 1698175906
transform -1 0 23072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__B1
timestamp 1698175906
transform 1 0 24192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__C1
timestamp 1698175906
transform -1 0 20048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__C2
timestamp 1698175906
transform -1 0 23520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0795__A1
timestamp 1698175906
transform 1 0 22400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__I
timestamp 1698175906
transform -1 0 27216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0799__A2
timestamp 1698175906
transform 1 0 23744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0800__I
timestamp 1698175906
transform 1 0 28224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0801__A1
timestamp 1698175906
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0802__B
timestamp 1698175906
transform 1 0 8064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0805__A2
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__A1
timestamp 1698175906
transform -1 0 11312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__B
timestamp 1698175906
transform -1 0 11760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0811__I
timestamp 1698175906
transform 1 0 23072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__A2
timestamp 1698175906
transform 1 0 24304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__A3
timestamp 1698175906
transform 1 0 25760 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0815__A2
timestamp 1698175906
transform 1 0 26880 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0816__A1
timestamp 1698175906
transform 1 0 25312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__A1
timestamp 1698175906
transform 1 0 16688 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__A2
timestamp 1698175906
transform 1 0 14784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__A1
timestamp 1698175906
transform 1 0 22400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__A2
timestamp 1698175906
transform 1 0 21952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0820__A1
timestamp 1698175906
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0820__A2
timestamp 1698175906
transform -1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__B
timestamp 1698175906
transform -1 0 17808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__C
timestamp 1698175906
transform -1 0 17360 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0826__A2
timestamp 1698175906
transform 1 0 19152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__A2
timestamp 1698175906
transform 1 0 16352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__B1
timestamp 1698175906
transform -1 0 17024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__A1
timestamp 1698175906
transform 1 0 10416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__C1
timestamp 1698175906
transform 1 0 19600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__C2
timestamp 1698175906
transform 1 0 21392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__I
timestamp 1698175906
transform 1 0 13664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__A1
timestamp 1698175906
transform 1 0 14448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__A1
timestamp 1698175906
transform -1 0 15232 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0837__I
timestamp 1698175906
transform 1 0 17472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__A2
timestamp 1698175906
transform 1 0 29008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__A1
timestamp 1698175906
transform 1 0 29232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__A2
timestamp 1698175906
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__A1
timestamp 1698175906
transform -1 0 12768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__A2
timestamp 1698175906
transform -1 0 21504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__B1
timestamp 1698175906
transform -1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__B2
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A1
timestamp 1698175906
transform -1 0 11648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A2
timestamp 1698175906
transform 1 0 11536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__A2
timestamp 1698175906
transform 1 0 29232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__A2
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__B2
timestamp 1698175906
transform 1 0 12992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A1
timestamp 1698175906
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A2
timestamp 1698175906
transform 1 0 21504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A1
timestamp 1698175906
transform 1 0 27552 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A2
timestamp 1698175906
transform 1 0 23744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__A1
timestamp 1698175906
transform 1 0 27104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__A2
timestamp 1698175906
transform 1 0 26656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__B
timestamp 1698175906
transform -1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__A1
timestamp 1698175906
transform 1 0 27216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__B1
timestamp 1698175906
transform 1 0 28784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__B2
timestamp 1698175906
transform 1 0 29232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A1
timestamp 1698175906
transform 1 0 29008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__B2
timestamp 1698175906
transform 1 0 7280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A1
timestamp 1698175906
transform -1 0 18144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__A1
timestamp 1698175906
transform 1 0 14560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__A2
timestamp 1698175906
transform 1 0 15008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__B1
timestamp 1698175906
transform 1 0 15456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__I
timestamp 1698175906
transform 1 0 15680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__A1
timestamp 1698175906
transform 1 0 21392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__I
timestamp 1698175906
transform 1 0 26880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A1
timestamp 1698175906
transform 1 0 18256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A2
timestamp 1698175906
transform 1 0 19264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__I
timestamp 1698175906
transform -1 0 22288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__A1
timestamp 1698175906
transform 1 0 17584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__I
timestamp 1698175906
transform -1 0 26656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__B1
timestamp 1698175906
transform 1 0 18480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__B2
timestamp 1698175906
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A2
timestamp 1698175906
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A1
timestamp 1698175906
transform -1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A2
timestamp 1698175906
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__A1
timestamp 1698175906
transform 1 0 28112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__A2
timestamp 1698175906
transform 1 0 28896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__B1
timestamp 1698175906
transform -1 0 17360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A2
timestamp 1698175906
transform 1 0 28112 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__B
timestamp 1698175906
transform 1 0 26992 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__A1
timestamp 1698175906
transform -1 0 7168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__A2
timestamp 1698175906
transform -1 0 6720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__A1
timestamp 1698175906
transform -1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__C1
timestamp 1698175906
transform -1 0 12656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__A2
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__A1
timestamp 1698175906
transform 1 0 16128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__A2
timestamp 1698175906
transform -1 0 14560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A1
timestamp 1698175906
transform 1 0 14896 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__B1
timestamp 1698175906
transform -1 0 15568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A2
timestamp 1698175906
transform 1 0 22848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A3
timestamp 1698175906
transform 1 0 22624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A4
timestamp 1698175906
transform 1 0 23072 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__A1
timestamp 1698175906
transform 1 0 24528 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A1
timestamp 1698175906
transform -1 0 24416 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A2
timestamp 1698175906
transform -1 0 23968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__A1
timestamp 1698175906
transform 1 0 24640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A2
timestamp 1698175906
transform -1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__A1
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A1
timestamp 1698175906
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A1
timestamp 1698175906
transform 1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A2
timestamp 1698175906
transform 1 0 24192 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__A1
timestamp 1698175906
transform 1 0 11088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__A2
timestamp 1698175906
transform 1 0 10080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A1
timestamp 1698175906
transform -1 0 8960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__B1
timestamp 1698175906
transform 1 0 11424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__B2
timestamp 1698175906
transform 1 0 12096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__A1
timestamp 1698175906
transform -1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__A2
timestamp 1698175906
transform 1 0 7056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__A2
timestamp 1698175906
transform 1 0 7504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__I
timestamp 1698175906
transform 1 0 14112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0938__I
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__A2
timestamp 1698175906
transform 1 0 10528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__B
timestamp 1698175906
transform 1 0 10080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A1
timestamp 1698175906
transform 1 0 10528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__B
timestamp 1698175906
transform 1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__A1
timestamp 1698175906
transform 1 0 4144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__A1
timestamp 1698175906
transform -1 0 4816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A3
timestamp 1698175906
transform 1 0 23072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__I
timestamp 1698175906
transform 1 0 30352 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__A2
timestamp 1698175906
transform 1 0 22624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__A1
timestamp 1698175906
transform 1 0 23184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__A2
timestamp 1698175906
transform 1 0 19936 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__A1
timestamp 1698175906
transform 1 0 19376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__B
timestamp 1698175906
transform 1 0 18032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0959__B2
timestamp 1698175906
transform 1 0 15008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0960__A1
timestamp 1698175906
transform 1 0 15456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A1
timestamp 1698175906
transform -1 0 3584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A3
timestamp 1698175906
transform 1 0 4592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A1
timestamp 1698175906
transform 1 0 29232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__A1
timestamp 1698175906
transform 1 0 28672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__A2
timestamp 1698175906
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__A2
timestamp 1698175906
transform 1 0 18816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__A1
timestamp 1698175906
transform 1 0 20272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__A2
timestamp 1698175906
transform -1 0 10752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A1
timestamp 1698175906
transform -1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A2
timestamp 1698175906
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__B1
timestamp 1698175906
transform -1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__A1
timestamp 1698175906
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__C2
timestamp 1698175906
transform 1 0 4592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__A4
timestamp 1698175906
transform 1 0 27104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A1
timestamp 1698175906
transform -1 0 17248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A1
timestamp 1698175906
transform -1 0 14224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A3
timestamp 1698175906
transform -1 0 20272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__A1
timestamp 1698175906
transform -1 0 16240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__B
timestamp 1698175906
transform -1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__A1
timestamp 1698175906
transform -1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__B1
timestamp 1698175906
transform 1 0 13664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__B2
timestamp 1698175906
transform -1 0 15008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0992__A1
timestamp 1698175906
transform -1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0994__A1
timestamp 1698175906
transform 1 0 22400 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A3
timestamp 1698175906
transform 1 0 22960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__A2
timestamp 1698175906
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__B
timestamp 1698175906
transform 1 0 28112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__C
timestamp 1698175906
transform 1 0 32144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__A1
timestamp 1698175906
transform -1 0 18928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__A3
timestamp 1698175906
transform 1 0 21840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A1
timestamp 1698175906
transform 1 0 18928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A2
timestamp 1698175906
transform -1 0 19600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__B2
timestamp 1698175906
transform 1 0 20832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1005__A1
timestamp 1698175906
transform -1 0 21168 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A1
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A1
timestamp 1698175906
transform -1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A3
timestamp 1698175906
transform -1 0 19824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A4
timestamp 1698175906
transform -1 0 18704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__C2
timestamp 1698175906
transform 1 0 23632 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1014__A3
timestamp 1698175906
transform 1 0 21504 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A1
timestamp 1698175906
transform -1 0 27888 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A1
timestamp 1698175906
transform 1 0 20496 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A1
timestamp 1698175906
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A1
timestamp 1698175906
transform 1 0 15344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__A1
timestamp 1698175906
transform 1 0 22512 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__I
timestamp 1698175906
transform 1 0 10416 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__I
timestamp 1698175906
transform 1 0 12768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__I
timestamp 1698175906
transform 1 0 12432 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A1
timestamp 1698175906
transform -1 0 12656 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A1
timestamp 1698175906
transform -1 0 12096 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1698175906
transform -1 0 11984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A1
timestamp 1698175906
transform 1 0 12768 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__A1
timestamp 1698175906
transform 1 0 11872 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A1
timestamp 1698175906
transform 1 0 11536 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I
timestamp 1698175906
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A1
timestamp 1698175906
transform -1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A1
timestamp 1698175906
transform 1 0 12320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__I
timestamp 1698175906
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__I
timestamp 1698175906
transform 1 0 34608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A1
timestamp 1698175906
transform 1 0 36288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698175906
transform 1 0 34720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698175906
transform -1 0 34160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__A1
timestamp 1698175906
transform -1 0 36848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__A1
timestamp 1698175906
transform 1 0 33936 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1061__A1
timestamp 1698175906
transform -1 0 36400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A2
timestamp 1698175906
transform 1 0 34048 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A1
timestamp 1698175906
transform 1 0 35392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__A2
timestamp 1698175906
transform -1 0 13440 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__I
timestamp 1698175906
transform 1 0 21728 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__I
timestamp 1698175906
transform 1 0 25760 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__I
timestamp 1698175906
transform 1 0 27440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__A1
timestamp 1698175906
transform 1 0 23408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698175906
transform 1 0 25536 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A1
timestamp 1698175906
transform 1 0 21952 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698175906
transform 1 0 27328 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__I
timestamp 1698175906
transform 1 0 38416 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__I
timestamp 1698175906
transform -1 0 38528 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__I
timestamp 1698175906
transform 1 0 38080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A1
timestamp 1698175906
transform 1 0 40320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A1
timestamp 1698175906
transform 1 0 40096 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__A1
timestamp 1698175906
transform 1 0 38640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A1
timestamp 1698175906
transform 1 0 40992 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__I
timestamp 1698175906
transform 1 0 29232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__I
timestamp 1698175906
transform 1 0 32592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__I
timestamp 1698175906
transform 1 0 37744 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A1
timestamp 1698175906
transform 1 0 28784 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A1
timestamp 1698175906
transform 1 0 29120 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__A1
timestamp 1698175906
transform 1 0 32480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__I
timestamp 1698175906
transform 1 0 37632 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A1
timestamp 1698175906
transform 1 0 32704 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__I
timestamp 1698175906
transform 1 0 38864 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__I
timestamp 1698175906
transform 1 0 38192 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A1
timestamp 1698175906
transform 1 0 38528 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1698175906
transform 1 0 40320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A1
timestamp 1698175906
transform 1 0 41216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__A1
timestamp 1698175906
transform 1 0 40320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__I
timestamp 1698175906
transform 1 0 15904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A1
timestamp 1698175906
transform 1 0 15344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__A1
timestamp 1698175906
transform 1 0 15344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1698175906
transform 1 0 18144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__A1
timestamp 1698175906
transform 1 0 19040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__I
timestamp 1698175906
transform 1 0 33040 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698175906
transform -1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1698175906
transform 1 0 36064 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__A1
timestamp 1698175906
transform 1 0 35616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__A1
timestamp 1698175906
transform 1 0 32144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__CLK
timestamp 1698175906
transform 1 0 5040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__CLK
timestamp 1698175906
transform 1 0 5040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__CLK
timestamp 1698175906
transform 1 0 8960 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__CLK
timestamp 1698175906
transform 1 0 39648 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__CLK
timestamp 1698175906
transform 1 0 33152 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__CLK
timestamp 1698175906
transform 1 0 36848 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__CLK
timestamp 1698175906
transform 1 0 36400 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__CLK
timestamp 1698175906
transform 1 0 36400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__CLK
timestamp 1698175906
transform 1 0 41664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__CLK
timestamp 1698175906
transform 1 0 40880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__CLK
timestamp 1698175906
transform 1 0 39872 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__CLK
timestamp 1698175906
transform 1 0 16800 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__CLK
timestamp 1698175906
transform 1 0 16464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__CLK
timestamp 1698175906
transform 1 0 21392 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__CLK
timestamp 1698175906
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__CLK
timestamp 1698175906
transform 1 0 37744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__CLK
timestamp 1698175906
transform 1 0 32368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 24192 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 27440 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 23072 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 33824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 7504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform -1 0 23184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform -1 0 25424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform -1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform -1 0 29904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform -1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform -1 0 34384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform -1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform -1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform -1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform -1 0 18704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform -1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform -1 0 11984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform -1 0 9744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform 1 0 1792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform 1 0 2464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698175906
transform 1 0 2464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698175906
transform 1 0 2464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698175906
transform 1 0 2464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698175906
transform 1 0 3136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698175906
transform -1 0 2240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698175906
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698175906
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698175906
transform 1 0 3136 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698175906
transform 1 0 1792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698175906
transform 1 0 2464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698175906
transform 1 0 1792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698175906
transform 1 0 1792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698175906
transform 1 0 2464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698175906
transform 1 0 2464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698175906
transform 1 0 2688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698175906
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698175906
transform 1 0 2464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698175906
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698175906
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698175906
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698175906
transform 1 0 3136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698175906
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698175906
transform 1 0 1792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698175906
transform 1 0 2464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698175906
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698175906
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698175906
transform -1 0 14224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698175906
transform -1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output49_I
timestamp 1698175906
transform -1 0 38976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1698175906
transform 1 0 43568 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1698175906
transform 1 0 45360 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698175906
transform -1 0 47824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1698175906
transform 1 0 50848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output54_I
timestamp 1698175906
transform 1 0 52080 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1698175906
transform -1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output56_I
timestamp 1698175906
transform 1 0 55216 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1698175906
transform -1 0 27216 0 1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1698175906
transform -1 0 22848 0 -1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1698175906
transform 1 0 33264 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1698175906
transform 1 0 33040 0 -1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_10 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_30 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698175906
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698175906
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698175906
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698175906
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698175906
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698175906
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1698175906
transform 1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_12
timestamp 1698175906
transform 1 0 2688 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_44
timestamp 1698175906
transform 1 0 6272 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_60
timestamp 1698175906
transform 1 0 8064 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_68
timestamp 1698175906
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698175906
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698175906
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698175906
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698175906
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698175906
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698175906
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6
timestamp 1698175906
transform 1 0 2016 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698175906
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698175906
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698175906
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698175906
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698175906
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698175906
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698175906
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698175906
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_10
timestamp 1698175906
transform 1 0 2464 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_42
timestamp 1698175906
transform 1 0 6048 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_58
timestamp 1698175906
transform 1 0 7840 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698175906
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698175906
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698175906
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698175906
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698175906
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698175906
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698175906
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698175906
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698175906
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698175906
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698175906
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698175906
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698175906
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698175906
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698175906
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698175906
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698175906
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698175906
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_12
timestamp 1698175906
transform 1 0 2688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698175906
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698175906
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698175906
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698175906
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698175906
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698175906
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698175906
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698175906
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698175906
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698175906
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698175906
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698175906
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698175906
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698175906
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698175906
transform 1 0 2688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698175906
transform 1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698175906
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698175906
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698175906
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698175906
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698175906
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698175906
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698175906
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698175906
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698175906
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698175906
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698175906
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698175906
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698175906
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698175906
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698175906
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698175906
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698175906
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698175906
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698175906
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_457
timestamp 1698175906
transform 1 0 52528 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_489
timestamp 1698175906
transform 1 0 56112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698175906
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698175906
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698175906
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698175906
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698175906
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698175906
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698175906
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698175906
transform 1 0 2688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698175906
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698175906
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698175906
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698175906
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698175906
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698175906
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698175906
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_505
timestamp 1698175906
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698175906
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698175906
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698175906
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698175906
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698175906
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698175906
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698175906
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698175906
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698175906
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_457
timestamp 1698175906
transform 1 0 52528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_489
timestamp 1698175906
transform 1 0 56112 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1698175906
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_8
timestamp 1698175906
transform 1 0 2240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_12
timestamp 1698175906
transform 1 0 2688 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_44
timestamp 1698175906
transform 1 0 6272 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_60
timestamp 1698175906
transform 1 0 8064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698175906
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698175906
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698175906
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698175906
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698175906
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698175906
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698175906
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698175906
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698175906
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698175906
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_457
timestamp 1698175906
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_489
timestamp 1698175906
transform 1 0 56112 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_505
timestamp 1698175906
transform 1 0 57904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_8
timestamp 1698175906
transform 1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_12
timestamp 1698175906
transform 1 0 2688 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_44
timestamp 1698175906
transform 1 0 6272 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698175906
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698175906
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698175906
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698175906
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698175906
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698175906
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698175906
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698175906
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698175906
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_457
timestamp 1698175906
transform 1 0 52528 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_489
timestamp 1698175906
transform 1 0 56112 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_505
timestamp 1698175906
transform 1 0 57904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698175906
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_12
timestamp 1698175906
transform 1 0 2688 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_44
timestamp 1698175906
transform 1 0 6272 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698175906
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698175906
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698175906
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698175906
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698175906
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698175906
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698175906
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698175906
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698175906
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_457
timestamp 1698175906
transform 1 0 52528 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_489
timestamp 1698175906
transform 1 0 56112 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_505
timestamp 1698175906
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698175906
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698175906
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698175906
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698175906
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698175906
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698175906
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698175906
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698175906
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698175906
transform 1 0 2688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698175906
transform 1 0 44016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698175906
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698175906
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_457
timestamp 1698175906
transform 1 0 52528 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_489
timestamp 1698175906
transform 1 0 56112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_505
timestamp 1698175906
transform 1 0 57904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698175906
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698175906
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698175906
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698175906
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698175906
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698175906
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_8
timestamp 1698175906
transform 1 0 2240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_12
timestamp 1698175906
transform 1 0 2688 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698175906
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698175906
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698175906
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_457
timestamp 1698175906
transform 1 0 52528 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_489
timestamp 1698175906
transform 1 0 56112 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_505
timestamp 1698175906
transform 1 0 57904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698175906
transform 1 0 14784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_124
timestamp 1698175906
transform 1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_133
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698175906
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_146
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_154
timestamp 1698175906
transform 1 0 18592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_161
timestamp 1698175906
transform 1 0 19376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_169
timestamp 1698175906
transform 1 0 20272 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_173
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_183
timestamp 1698175906
transform 1 0 21840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_187
timestamp 1698175906
transform 1 0 22288 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_191
timestamp 1698175906
transform 1 0 22736 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_194
timestamp 1698175906
transform 1 0 23072 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698175906
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698175906
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698175906
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698175906
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698175906
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698175906
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698175906
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698175906
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_85
timestamp 1698175906
transform 1 0 10864 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_89
timestamp 1698175906
transform 1 0 11312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_93
timestamp 1698175906
transform 1 0 11760 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_129
timestamp 1698175906
transform 1 0 15792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_192
timestamp 1698175906
transform 1 0 22848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_194
timestamp 1698175906
transform 1 0 23072 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_215
timestamp 1698175906
transform 1 0 25424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_219
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_235
timestamp 1698175906
transform 1 0 27664 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698175906
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698175906
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698175906
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_457
timestamp 1698175906
transform 1 0 52528 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_489
timestamp 1698175906
transform 1 0 56112 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_505
timestamp 1698175906
transform 1 0 57904 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698175906
transform 1 0 10976 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_89
timestamp 1698175906
transform 1 0 11312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_220
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_224
timestamp 1698175906
transform 1 0 26432 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_256
timestamp 1698175906
transform 1 0 30016 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_272
timestamp 1698175906
transform 1 0 31808 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698175906
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698175906
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698175906
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698175906
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698175906
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698175906
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698175906
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698175906
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698175906
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_59
timestamp 1698175906
transform 1 0 7952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698175906
transform 1 0 13552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_118
timestamp 1698175906
transform 1 0 14560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_159
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_228
timestamp 1698175906
transform 1 0 26880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_232
timestamp 1698175906
transform 1 0 27328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_234
timestamp 1698175906
transform 1 0 27552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_251
timestamp 1698175906
transform 1 0 29456 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698175906
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698175906
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698175906
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_457
timestamp 1698175906
transform 1 0 52528 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_489
timestamp 1698175906
transform 1 0 56112 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_505
timestamp 1698175906
transform 1 0 57904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_34
timestamp 1698175906
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_44
timestamp 1698175906
transform 1 0 6272 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_48
timestamp 1698175906
transform 1 0 6720 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_80
timestamp 1698175906
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_84
timestamp 1698175906
transform 1 0 10752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_112
timestamp 1698175906
transform 1 0 13888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_116
timestamp 1698175906
transform 1 0 14336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_120
timestamp 1698175906
transform 1 0 14784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698175906
transform 1 0 16240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_137
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_151
timestamp 1698175906
transform 1 0 18256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_155
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_157
timestamp 1698175906
transform 1 0 18928 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_160
timestamp 1698175906
transform 1 0 19264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_164
timestamp 1698175906
transform 1 0 19712 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_168
timestamp 1698175906
transform 1 0 20160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_172
timestamp 1698175906
transform 1 0 20608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_184
timestamp 1698175906
transform 1 0 21952 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_193
timestamp 1698175906
transform 1 0 22960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_197
timestamp 1698175906
transform 1 0 23408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_205
timestamp 1698175906
transform 1 0 24304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_222
timestamp 1698175906
transform 1 0 26208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_226
timestamp 1698175906
transform 1 0 26656 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_258
timestamp 1698175906
transform 1 0 30240 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_274
timestamp 1698175906
transform 1 0 32032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698175906
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698175906
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698175906
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698175906
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698175906
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698175906
transform 1 0 56448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698175906
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_27
timestamp 1698175906
transform 1 0 4368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_31
timestamp 1698175906
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_47
timestamp 1698175906
transform 1 0 6608 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_55
timestamp 1698175906
transform 1 0 7504 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_59
timestamp 1698175906
transform 1 0 7952 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_62
timestamp 1698175906
transform 1 0 8288 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_76
timestamp 1698175906
transform 1 0 9856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_80
timestamp 1698175906
transform 1 0 10304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_84
timestamp 1698175906
transform 1 0 10752 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_92
timestamp 1698175906
transform 1 0 11648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_94
timestamp 1698175906
transform 1 0 11872 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698175906
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_115
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_132
timestamp 1698175906
transform 1 0 16128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_138
timestamp 1698175906
transform 1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_142
timestamp 1698175906
transform 1 0 17248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_144
timestamp 1698175906
transform 1 0 17472 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_147
timestamp 1698175906
transform 1 0 17808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_159
timestamp 1698175906
transform 1 0 19152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_163
timestamp 1698175906
transform 1 0 19600 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698175906
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698175906
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698175906
transform 1 0 21840 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_186
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_194
timestamp 1698175906
transform 1 0 23072 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_198
timestamp 1698175906
transform 1 0 23520 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_223
timestamp 1698175906
transform 1 0 26320 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_227
timestamp 1698175906
transform 1 0 26768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_231
timestamp 1698175906
transform 1 0 27216 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698175906
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698175906
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698175906
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_457
timestamp 1698175906
transform 1 0 52528 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_489
timestamp 1698175906
transform 1 0 56112 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_505
timestamp 1698175906
transform 1 0 57904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_8
timestamp 1698175906
transform 1 0 2240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_12
timestamp 1698175906
transform 1 0 2688 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_20
timestamp 1698175906
transform 1 0 3584 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_24
timestamp 1698175906
transform 1 0 4032 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_27
timestamp 1698175906
transform 1 0 4368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_54
timestamp 1698175906
transform 1 0 7392 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_86
timestamp 1698175906
transform 1 0 10976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_92
timestamp 1698175906
transform 1 0 11648 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_182
timestamp 1698175906
transform 1 0 21728 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_190
timestamp 1698175906
transform 1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_194
timestamp 1698175906
transform 1 0 23072 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_202
timestamp 1698175906
transform 1 0 23968 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_221
timestamp 1698175906
transform 1 0 26096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_237
timestamp 1698175906
transform 1 0 27888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_241
timestamp 1698175906
transform 1 0 28336 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_265
timestamp 1698175906
transform 1 0 31024 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_273
timestamp 1698175906
transform 1 0 31920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698175906
transform 1 0 32368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698175906
transform 1 0 40768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698175906
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698175906
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698175906
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_492
timestamp 1698175906
transform 1 0 56448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698175906
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_6
timestamp 1698175906
transform 1 0 2016 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_25
timestamp 1698175906
transform 1 0 4144 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_33
timestamp 1698175906
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_41
timestamp 1698175906
transform 1 0 5936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_90
timestamp 1698175906
transform 1 0 11424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_94
timestamp 1698175906
transform 1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_98
timestamp 1698175906
transform 1 0 12320 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_100
timestamp 1698175906
transform 1 0 12544 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698175906
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_115
timestamp 1698175906
transform 1 0 14224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_127
timestamp 1698175906
transform 1 0 15568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_129
timestamp 1698175906
transform 1 0 15792 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_138
timestamp 1698175906
transform 1 0 16800 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_146
timestamp 1698175906
transform 1 0 17696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_150
timestamp 1698175906
transform 1 0 18144 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_158
timestamp 1698175906
transform 1 0 19040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_162
timestamp 1698175906
transform 1 0 19488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_166
timestamp 1698175906
transform 1 0 19936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_191
timestamp 1698175906
transform 1 0 22736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_193
timestamp 1698175906
transform 1 0 22960 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_210
timestamp 1698175906
transform 1 0 24864 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_214
timestamp 1698175906
transform 1 0 25312 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_226
timestamp 1698175906
transform 1 0 26656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_230
timestamp 1698175906
transform 1 0 27104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_232
timestamp 1698175906
transform 1 0 27328 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_235
timestamp 1698175906
transform 1 0 27664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698175906
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_260
timestamp 1698175906
transform 1 0 30464 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_292
timestamp 1698175906
transform 1 0 34048 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_308
timestamp 1698175906
transform 1 0 35840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698175906
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698175906
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698175906
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698175906
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698175906
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_457
timestamp 1698175906
transform 1 0 52528 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_489
timestamp 1698175906
transform 1 0 56112 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_505
timestamp 1698175906
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_6
timestamp 1698175906
transform 1 0 2016 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_47
timestamp 1698175906
transform 1 0 6608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698175906
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_88
timestamp 1698175906
transform 1 0 11200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_90
timestamp 1698175906
transform 1 0 11424 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_101
timestamp 1698175906
transform 1 0 12656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_114
timestamp 1698175906
transform 1 0 14112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_125
timestamp 1698175906
transform 1 0 15344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_127
timestamp 1698175906
transform 1 0 15568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_130
timestamp 1698175906
transform 1 0 15904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_134
timestamp 1698175906
transform 1 0 16352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_138
timestamp 1698175906
transform 1 0 16800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_150
timestamp 1698175906
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_154
timestamp 1698175906
transform 1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_156
timestamp 1698175906
transform 1 0 18816 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_159
timestamp 1698175906
transform 1 0 19152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_172
timestamp 1698175906
transform 1 0 20608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_184
timestamp 1698175906
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_188
timestamp 1698175906
transform 1 0 22400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_192
timestamp 1698175906
transform 1 0 22848 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_198
timestamp 1698175906
transform 1 0 23520 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_207
timestamp 1698175906
transform 1 0 24528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698175906
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_218
timestamp 1698175906
transform 1 0 25760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_222
timestamp 1698175906
transform 1 0 26208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_228
timestamp 1698175906
transform 1 0 26880 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_256
timestamp 1698175906
transform 1 0 30016 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_272
timestamp 1698175906
transform 1 0 31808 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_290
timestamp 1698175906
transform 1 0 33824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_329
timestamp 1698175906
transform 1 0 38192 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_345
timestamp 1698175906
transform 1 0 39984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698175906
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698175906
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698175906
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698175906
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698175906
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698175906
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698175906
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_14
timestamp 1698175906
transform 1 0 2912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_18
timestamp 1698175906
transform 1 0 3360 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_22
timestamp 1698175906
transform 1 0 3808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_26
timestamp 1698175906
transform 1 0 4256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_39
timestamp 1698175906
transform 1 0 5712 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_51
timestamp 1698175906
transform 1 0 7056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_53
timestamp 1698175906
transform 1 0 7280 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_79
timestamp 1698175906
transform 1 0 10192 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_85
timestamp 1698175906
transform 1 0 10864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_98
timestamp 1698175906
transform 1 0 12320 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698175906
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_115
timestamp 1698175906
transform 1 0 14224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_119
timestamp 1698175906
transform 1 0 14672 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_123
timestamp 1698175906
transform 1 0 15120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_127
timestamp 1698175906
transform 1 0 15568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_135
timestamp 1698175906
transform 1 0 16464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_139
timestamp 1698175906
transform 1 0 16912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_186
timestamp 1698175906
transform 1 0 22176 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_227
timestamp 1698175906
transform 1 0 26768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_231
timestamp 1698175906
transform 1 0 27216 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_251
timestamp 1698175906
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_253
timestamp 1698175906
transform 1 0 29680 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_276
timestamp 1698175906
transform 1 0 32256 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_292
timestamp 1698175906
transform 1 0 34048 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_302
timestamp 1698175906
transform 1 0 35168 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_306
timestamp 1698175906
transform 1 0 35616 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1698175906
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698175906
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698175906
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698175906
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_457
timestamp 1698175906
transform 1 0 52528 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_489
timestamp 1698175906
transform 1 0 56112 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_505
timestamp 1698175906
transform 1 0 57904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_4
timestamp 1698175906
transform 1 0 1792 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_53
timestamp 1698175906
transform 1 0 7280 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_57
timestamp 1698175906
transform 1 0 7728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_61
timestamp 1698175906
transform 1 0 8176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_63
timestamp 1698175906
transform 1 0 8400 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_104
timestamp 1698175906
transform 1 0 12992 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_108
timestamp 1698175906
transform 1 0 13440 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_120
timestamp 1698175906
transform 1 0 14784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_124
timestamp 1698175906
transform 1 0 15232 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_128
timestamp 1698175906
transform 1 0 15680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_130
timestamp 1698175906
transform 1 0 15904 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_151
timestamp 1698175906
transform 1 0 18256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_161
timestamp 1698175906
transform 1 0 19376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_165
timestamp 1698175906
transform 1 0 19824 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_177
timestamp 1698175906
transform 1 0 21168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_181
timestamp 1698175906
transform 1 0 21616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_185
timestamp 1698175906
transform 1 0 22064 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_201
timestamp 1698175906
transform 1 0 23856 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_203
timestamp 1698175906
transform 1 0 24080 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_228
timestamp 1698175906
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_230
timestamp 1698175906
transform 1 0 27104 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_239
timestamp 1698175906
transform 1 0 28112 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_241
timestamp 1698175906
transform 1 0 28336 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_252
timestamp 1698175906
transform 1 0 29568 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_268
timestamp 1698175906
transform 1 0 31360 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_333
timestamp 1698175906
transform 1 0 38640 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698175906
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698175906
transform 1 0 40768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698175906
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698175906
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698175906
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698175906
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698175906
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_6
timestamp 1698175906
transform 1 0 2016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_8
timestamp 1698175906
transform 1 0 2240 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_25
timestamp 1698175906
transform 1 0 4144 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698175906
transform 1 0 5040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_53
timestamp 1698175906
transform 1 0 7280 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_57
timestamp 1698175906
transform 1 0 7728 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698175906
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_126
timestamp 1698175906
transform 1 0 15456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_160
timestamp 1698175906
transform 1 0 19264 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_181
timestamp 1698175906
transform 1 0 21616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_185
timestamp 1698175906
transform 1 0 22064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_195
timestamp 1698175906
transform 1 0 23184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_197
timestamp 1698175906
transform 1 0 23408 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698175906
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_255
timestamp 1698175906
transform 1 0 29904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_257
timestamp 1698175906
transform 1 0 30128 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_266
timestamp 1698175906
transform 1 0 31136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_274
timestamp 1698175906
transform 1 0 32032 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698175906
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698175906
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_354
timestamp 1698175906
transform 1 0 40992 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_370
timestamp 1698175906
transform 1 0 42784 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_378
timestamp 1698175906
transform 1 0 43680 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698175906
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698175906
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698175906
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698175906
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_457
timestamp 1698175906
transform 1 0 52528 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_489
timestamp 1698175906
transform 1 0 56112 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_505
timestamp 1698175906
transform 1 0 57904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_51
timestamp 1698175906
transform 1 0 7056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_55
timestamp 1698175906
transform 1 0 7504 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_59
timestamp 1698175906
transform 1 0 7952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_61
timestamp 1698175906
transform 1 0 8176 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_76
timestamp 1698175906
transform 1 0 9856 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_110
timestamp 1698175906
transform 1 0 13664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_112
timestamp 1698175906
transform 1 0 13888 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_123
timestamp 1698175906
transform 1 0 15120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_127
timestamp 1698175906
transform 1 0 15568 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_131
timestamp 1698175906
transform 1 0 16016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_133
timestamp 1698175906
transform 1 0 16240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_157
timestamp 1698175906
transform 1 0 18928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_161
timestamp 1698175906
transform 1 0 19376 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_177
timestamp 1698175906
transform 1 0 21168 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_203
timestamp 1698175906
transform 1 0 24080 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_207
timestamp 1698175906
transform 1 0 24528 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_244
timestamp 1698175906
transform 1 0 28672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_248
timestamp 1698175906
transform 1 0 29120 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_319
timestamp 1698175906
transform 1 0 37072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698175906
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_352
timestamp 1698175906
transform 1 0 40768 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698175906
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698175906
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698175906
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698175906
transform 1 0 56448 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698175906
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698175906
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_39
timestamp 1698175906
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_72
timestamp 1698175906
transform 1 0 9408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_76
timestamp 1698175906
transform 1 0 9856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_80
timestamp 1698175906
transform 1 0 10304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_88
timestamp 1698175906
transform 1 0 11200 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_92
timestamp 1698175906
transform 1 0 11648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_94
timestamp 1698175906
transform 1 0 11872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_97
timestamp 1698175906
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_109
timestamp 1698175906
transform 1 0 13552 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_112
timestamp 1698175906
transform 1 0 13888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_116
timestamp 1698175906
transform 1 0 14336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_120
timestamp 1698175906
transform 1 0 14784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_124
timestamp 1698175906
transform 1 0 15232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_128
timestamp 1698175906
transform 1 0 15680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_132
timestamp 1698175906
transform 1 0 16128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_136
timestamp 1698175906
transform 1 0 16576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_138
timestamp 1698175906
transform 1 0 16800 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_160
timestamp 1698175906
transform 1 0 19264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_164
timestamp 1698175906
transform 1 0 19712 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_168
timestamp 1698175906
transform 1 0 20160 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_179
timestamp 1698175906
transform 1 0 21392 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_182
timestamp 1698175906
transform 1 0 21728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_186
timestamp 1698175906
transform 1 0 22176 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_230
timestamp 1698175906
transform 1 0 27104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_232
timestamp 1698175906
transform 1 0 27328 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698175906
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698175906
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_251
timestamp 1698175906
transform 1 0 29456 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698175906
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_257
timestamp 1698175906
transform 1 0 30128 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_266
timestamp 1698175906
transform 1 0 31136 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_274
timestamp 1698175906
transform 1 0 32032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_292
timestamp 1698175906
transform 1 0 34048 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_296
timestamp 1698175906
transform 1 0 34496 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_359
timestamp 1698175906
transform 1 0 41552 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_375
timestamp 1698175906
transform 1 0 43344 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1698175906
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698175906
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698175906
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_457
timestamp 1698175906
transform 1 0 52528 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_489
timestamp 1698175906
transform 1 0 56112 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_505
timestamp 1698175906
transform 1 0 57904 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_8
timestamp 1698175906
transform 1 0 2240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_12
timestamp 1698175906
transform 1 0 2688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_16
timestamp 1698175906
transform 1 0 3136 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_25
timestamp 1698175906
transform 1 0 4144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_33
timestamp 1698175906
transform 1 0 5040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_43
timestamp 1698175906
transform 1 0 6160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_45
timestamp 1698175906
transform 1 0 6384 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_48
timestamp 1698175906
transform 1 0 6720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_60
timestamp 1698175906
transform 1 0 8064 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698175906
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_85
timestamp 1698175906
transform 1 0 10864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_89
timestamp 1698175906
transform 1 0 11312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_101
timestamp 1698175906
transform 1 0 12656 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_134
timestamp 1698175906
transform 1 0 16352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698175906
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_147
timestamp 1698175906
transform 1 0 17808 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_159
timestamp 1698175906
transform 1 0 19152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_161
timestamp 1698175906
transform 1 0 19376 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_205
timestamp 1698175906
transform 1 0 24304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_207
timestamp 1698175906
transform 1 0 24528 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_227
timestamp 1698175906
transform 1 0 26768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_243
timestamp 1698175906
transform 1 0 28560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_247
timestamp 1698175906
transform 1 0 29008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_251
timestamp 1698175906
transform 1 0 29456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_253
timestamp 1698175906
transform 1 0 29680 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_270
timestamp 1698175906
transform 1 0 31584 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_322
timestamp 1698175906
transform 1 0 37408 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_345
timestamp 1698175906
transform 1 0 39984 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698175906
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698175906
transform 1 0 40768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698175906
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698175906
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698175906
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698175906
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698175906
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_6
timestamp 1698175906
transform 1 0 2016 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_16
timestamp 1698175906
transform 1 0 3136 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698175906
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_67
timestamp 1698175906
transform 1 0 8848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_93
timestamp 1698175906
transform 1 0 11760 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_164
timestamp 1698175906
transform 1 0 19712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_166
timestamp 1698175906
transform 1 0 19936 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_179
timestamp 1698175906
transform 1 0 21392 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_252
timestamp 1698175906
transform 1 0 29568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_266
timestamp 1698175906
transform 1 0 31136 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_268
timestamp 1698175906
transform 1 0 31360 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698175906
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_319
timestamp 1698175906
transform 1 0 37072 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_365
timestamp 1698175906
transform 1 0 42224 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_381
timestamp 1698175906
transform 1 0 44016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698175906
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698175906
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_457
timestamp 1698175906
transform 1 0 52528 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_489
timestamp 1698175906
transform 1 0 56112 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_505
timestamp 1698175906
transform 1 0 57904 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_6
timestamp 1698175906
transform 1 0 2016 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_23
timestamp 1698175906
transform 1 0 3920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_27
timestamp 1698175906
transform 1 0 4368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_31
timestamp 1698175906
transform 1 0 4816 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_35
timestamp 1698175906
transform 1 0 5264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_37
timestamp 1698175906
transform 1 0 5488 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_46
timestamp 1698175906
transform 1 0 6496 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_54
timestamp 1698175906
transform 1 0 7392 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_63
timestamp 1698175906
transform 1 0 8400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_67
timestamp 1698175906
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698175906
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_81
timestamp 1698175906
transform 1 0 10416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_85
timestamp 1698175906
transform 1 0 10864 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_89
timestamp 1698175906
transform 1 0 11312 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_92
timestamp 1698175906
transform 1 0 11648 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_98
timestamp 1698175906
transform 1 0 12320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_102
timestamp 1698175906
transform 1 0 12768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_106
timestamp 1698175906
transform 1 0 13216 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_123
timestamp 1698175906
transform 1 0 15120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_127
timestamp 1698175906
transform 1 0 15568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_135
timestamp 1698175906
transform 1 0 16464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698175906
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_162
timestamp 1698175906
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_221
timestamp 1698175906
transform 1 0 26096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_225
timestamp 1698175906
transform 1 0 26544 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_228
timestamp 1698175906
transform 1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_238
timestamp 1698175906
transform 1 0 28000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_242
timestamp 1698175906
transform 1 0 28448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_246
timestamp 1698175906
transform 1 0 28896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_250
timestamp 1698175906
transform 1 0 29344 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_266
timestamp 1698175906
transform 1 0 31136 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_274
timestamp 1698175906
transform 1 0 32032 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_278
timestamp 1698175906
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_352
timestamp 1698175906
transform 1 0 40768 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698175906
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698175906
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698175906
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698175906
transform 1 0 56448 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698175906
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_29
timestamp 1698175906
transform 1 0 4592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_33
timestamp 1698175906
transform 1 0 5040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_43
timestamp 1698175906
transform 1 0 6160 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_66
timestamp 1698175906
transform 1 0 8736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_70
timestamp 1698175906
transform 1 0 9184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_78
timestamp 1698175906
transform 1 0 10080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_80
timestamp 1698175906
transform 1 0 10304 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_83
timestamp 1698175906
transform 1 0 10640 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_99
timestamp 1698175906
transform 1 0 12432 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_109
timestamp 1698175906
transform 1 0 13552 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_117
timestamp 1698175906
transform 1 0 14448 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_133
timestamp 1698175906
transform 1 0 16240 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_141
timestamp 1698175906
transform 1 0 17136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_143
timestamp 1698175906
transform 1 0 17360 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_153
timestamp 1698175906
transform 1 0 18480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_155
timestamp 1698175906
transform 1 0 18704 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_158
timestamp 1698175906
transform 1 0 19040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_162
timestamp 1698175906
transform 1 0 19488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_166
timestamp 1698175906
transform 1 0 19936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_181
timestamp 1698175906
transform 1 0 21616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_232
timestamp 1698175906
transform 1 0 27328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698175906
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_251
timestamp 1698175906
transform 1 0 29456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_255
timestamp 1698175906
transform 1 0 29904 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_263
timestamp 1698175906
transform 1 0 30800 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_267
timestamp 1698175906
transform 1 0 31248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_269
timestamp 1698175906
transform 1 0 31472 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_278
timestamp 1698175906
transform 1 0 32480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_288
timestamp 1698175906
transform 1 0 33600 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_325
timestamp 1698175906
transform 1 0 37744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_343
timestamp 1698175906
transform 1 0 39760 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_375
timestamp 1698175906
transform 1 0 43344 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_383
timestamp 1698175906
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698175906
transform 1 0 44688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698175906
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_457
timestamp 1698175906
transform 1 0 52528 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_489
timestamp 1698175906
transform 1 0 56112 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_505
timestamp 1698175906
transform 1 0 57904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_8
timestamp 1698175906
transform 1 0 2240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_14
timestamp 1698175906
transform 1 0 2912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_18
timestamp 1698175906
transform 1 0 3360 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_34
timestamp 1698175906
transform 1 0 5152 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_42
timestamp 1698175906
transform 1 0 6048 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_45
timestamp 1698175906
transform 1 0 6384 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_49
timestamp 1698175906
transform 1 0 6832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_51
timestamp 1698175906
transform 1 0 7056 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_83
timestamp 1698175906
transform 1 0 10640 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_91
timestamp 1698175906
transform 1 0 11536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_98
timestamp 1698175906
transform 1 0 12320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_102
timestamp 1698175906
transform 1 0 12768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_106
timestamp 1698175906
transform 1 0 13216 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_114
timestamp 1698175906
transform 1 0 14112 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_118
timestamp 1698175906
transform 1 0 14560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698175906
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698175906
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_155
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 25536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_290
timestamp 1698175906
transform 1 0 33824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_292
timestamp 1698175906
transform 1 0 34048 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_332
timestamp 1698175906
transform 1 0 38528 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698175906
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698175906
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698175906
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698175906
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698175906
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698175906
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_8
timestamp 1698175906
transform 1 0 2240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_33
timestamp 1698175906
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_62
timestamp 1698175906
transform 1 0 8288 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_80
timestamp 1698175906
transform 1 0 10304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_100
timestamp 1698175906
transform 1 0 12544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_132
timestamp 1698175906
transform 1 0 16128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_136
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_149
timestamp 1698175906
transform 1 0 18032 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_160
timestamp 1698175906
transform 1 0 19264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698175906
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_177
timestamp 1698175906
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_181
timestamp 1698175906
transform 1 0 21616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_185
timestamp 1698175906
transform 1 0 22064 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_187
timestamp 1698175906
transform 1 0 22288 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_190
timestamp 1698175906
transform 1 0 22624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_194
timestamp 1698175906
transform 1 0 23072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_198
timestamp 1698175906
transform 1 0 23520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698175906
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_251
timestamp 1698175906
transform 1 0 29456 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698175906
transform 1 0 30800 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698175906
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_277
timestamp 1698175906
transform 1 0 32368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_297
timestamp 1698175906
transform 1 0 34608 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698175906
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_317
timestamp 1698175906
transform 1 0 36848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_333
timestamp 1698175906
transform 1 0 38640 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_365
timestamp 1698175906
transform 1 0 42224 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698175906
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698175906
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698175906
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_457
timestamp 1698175906
transform 1 0 52528 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_489
timestamp 1698175906
transform 1 0 56112 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_505
timestamp 1698175906
transform 1 0 57904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_2
timestamp 1698175906
transform 1 0 1568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_6
timestamp 1698175906
transform 1 0 2016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_14
timestamp 1698175906
transform 1 0 2912 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_24
timestamp 1698175906
transform 1 0 4032 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_28
timestamp 1698175906
transform 1 0 4480 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_32
timestamp 1698175906
transform 1 0 4928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_62
timestamp 1698175906
transform 1 0 8288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698175906
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_72
timestamp 1698175906
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_88
timestamp 1698175906
transform 1 0 11200 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_106
timestamp 1698175906
transform 1 0 13216 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_110
timestamp 1698175906
transform 1 0 13664 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_128
timestamp 1698175906
transform 1 0 15680 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698175906
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698175906
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_146
timestamp 1698175906
transform 1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_150
timestamp 1698175906
transform 1 0 18144 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_154
timestamp 1698175906
transform 1 0 18592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_157
timestamp 1698175906
transform 1 0 18928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_163
timestamp 1698175906
transform 1 0 19600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_167
timestamp 1698175906
transform 1 0 20048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_171
timestamp 1698175906
transform 1 0 20496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_173
timestamp 1698175906
transform 1 0 20720 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_193
timestamp 1698175906
transform 1 0 22960 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_202
timestamp 1698175906
transform 1 0 23968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_206
timestamp 1698175906
transform 1 0 24416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_235
timestamp 1698175906
transform 1 0 27664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_245
timestamp 1698175906
transform 1 0 28784 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_249
timestamp 1698175906
transform 1 0 29232 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_253
timestamp 1698175906
transform 1 0 29680 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_261
timestamp 1698175906
transform 1 0 30576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_263
timestamp 1698175906
transform 1 0 30800 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_282
timestamp 1698175906
transform 1 0 32928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_286
timestamp 1698175906
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_320
timestamp 1698175906
transform 1 0 37184 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698175906
transform 1 0 40768 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698175906
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698175906
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698175906
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698175906
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698175906
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_2
timestamp 1698175906
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_10
timestamp 1698175906
transform 1 0 2464 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_37
timestamp 1698175906
transform 1 0 5488 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_41
timestamp 1698175906
transform 1 0 5936 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_76
timestamp 1698175906
transform 1 0 9856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_92
timestamp 1698175906
transform 1 0 11648 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_102
timestamp 1698175906
transform 1 0 12768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698175906
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698175906
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1698175906
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_113
timestamp 1698175906
transform 1 0 14000 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_116
timestamp 1698175906
transform 1 0 14336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_160
timestamp 1698175906
transform 1 0 19264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_164
timestamp 1698175906
transform 1 0 19712 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_172
timestamp 1698175906
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698175906
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_191
timestamp 1698175906
transform 1 0 22736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_232
timestamp 1698175906
transform 1 0 27328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_234
timestamp 1698175906
transform 1 0 27552 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_247
timestamp 1698175906
transform 1 0 29008 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_308
timestamp 1698175906
transform 1 0 35840 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1698175906
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698175906
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698175906
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698175906
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698175906
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698175906
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_457
timestamp 1698175906
transform 1 0 52528 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_489
timestamp 1698175906
transform 1 0 56112 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_505
timestamp 1698175906
transform 1 0 57904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_8
timestamp 1698175906
transform 1 0 2240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_12
timestamp 1698175906
transform 1 0 2688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_16
timestamp 1698175906
transform 1 0 3136 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_72
timestamp 1698175906
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_110
timestamp 1698175906
transform 1 0 13664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_122
timestamp 1698175906
transform 1 0 15008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698175906
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_148
timestamp 1698175906
transform 1 0 17920 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_163
timestamp 1698175906
transform 1 0 19600 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_171
timestamp 1698175906
transform 1 0 20496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_177
timestamp 1698175906
transform 1 0 21168 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_185
timestamp 1698175906
transform 1 0 22064 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_189
timestamp 1698175906
transform 1 0 22512 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_192
timestamp 1698175906
transform 1 0 22848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_196
timestamp 1698175906
transform 1 0 23296 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_200
timestamp 1698175906
transform 1 0 23744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_204
timestamp 1698175906
transform 1 0 24192 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698175906
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_228
timestamp 1698175906
transform 1 0 26880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_232
timestamp 1698175906
transform 1 0 27328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_234
timestamp 1698175906
transform 1 0 27552 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698175906
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_290
timestamp 1698175906
transform 1 0 33824 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_309
timestamp 1698175906
transform 1 0 35952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_313
timestamp 1698175906
transform 1 0 36400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_317
timestamp 1698175906
transform 1 0 36848 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698175906
transform 1 0 40432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698175906
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698175906
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698175906
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698175906
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698175906
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698175906
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_14
timestamp 1698175906
transform 1 0 2912 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_30
timestamp 1698175906
transform 1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698175906
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698175906
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_79
timestamp 1698175906
transform 1 0 10192 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_87
timestamp 1698175906
transform 1 0 11088 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_91
timestamp 1698175906
transform 1 0 11536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_102
timestamp 1698175906
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698175906
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698175906
transform 1 0 13328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_121
timestamp 1698175906
transform 1 0 14896 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_125
timestamp 1698175906
transform 1 0 15344 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_168
timestamp 1698175906
transform 1 0 20160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_187
timestamp 1698175906
transform 1 0 22288 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_191
timestamp 1698175906
transform 1 0 22736 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_226
timestamp 1698175906
transform 1 0 26656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_230
timestamp 1698175906
transform 1 0 27104 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_233
timestamp 1698175906
transform 1 0 27440 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_237
timestamp 1698175906
transform 1 0 27888 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_241
timestamp 1698175906
transform 1 0 28336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_297
timestamp 1698175906
transform 1 0 34608 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698175906
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_346
timestamp 1698175906
transform 1 0 40096 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_378
timestamp 1698175906
transform 1 0 43680 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_382
timestamp 1698175906
transform 1 0 44128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698175906
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698175906
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698175906
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_457
timestamp 1698175906
transform 1 0 52528 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_489
timestamp 1698175906
transform 1 0 56112 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_505
timestamp 1698175906
transform 1 0 57904 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_2
timestamp 1698175906
transform 1 0 1568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_6
timestamp 1698175906
transform 1 0 2016 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_16
timestamp 1698175906
transform 1 0 3136 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_26
timestamp 1698175906
transform 1 0 4256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_30
timestamp 1698175906
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_32
timestamp 1698175906
transform 1 0 4928 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_72
timestamp 1698175906
transform 1 0 9408 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_80
timestamp 1698175906
transform 1 0 10304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_113
timestamp 1698175906
transform 1 0 14000 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_129
timestamp 1698175906
transform 1 0 15792 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_133
timestamp 1698175906
transform 1 0 16240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_142
timestamp 1698175906
transform 1 0 17248 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_159
timestamp 1698175906
transform 1 0 19152 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_163
timestamp 1698175906
transform 1 0 19600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_165
timestamp 1698175906
transform 1 0 19824 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_177
timestamp 1698175906
transform 1 0 21168 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_179
timestamp 1698175906
transform 1 0 21392 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_193
timestamp 1698175906
transform 1 0 22960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_197
timestamp 1698175906
transform 1 0 23408 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_205
timestamp 1698175906
transform 1 0 24304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_207
timestamp 1698175906
transform 1 0 24528 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_212
timestamp 1698175906
transform 1 0 25088 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_226
timestamp 1698175906
transform 1 0 26656 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_230
timestamp 1698175906
transform 1 0 27104 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_273
timestamp 1698175906
transform 1 0 31920 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_277
timestamp 1698175906
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698175906
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698175906
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_286
timestamp 1698175906
transform 1 0 33376 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_290
timestamp 1698175906
transform 1 0 33824 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_299
timestamp 1698175906
transform 1 0 34832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_310
timestamp 1698175906
transform 1 0 36064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_314
timestamp 1698175906
transform 1 0 36512 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_330
timestamp 1698175906
transform 1 0 38304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_338
timestamp 1698175906
transform 1 0 39200 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_342
timestamp 1698175906
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698175906
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_381
timestamp 1698175906
transform 1 0 44016 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_413
timestamp 1698175906
transform 1 0 47600 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_417
timestamp 1698175906
transform 1 0 48048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698175906
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_422
timestamp 1698175906
transform 1 0 48608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_486
timestamp 1698175906
transform 1 0 55776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698175906
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698175906
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_8
timestamp 1698175906
transform 1 0 2240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_10
timestamp 1698175906
transform 1 0 2464 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_16
timestamp 1698175906
transform 1 0 3136 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_32
timestamp 1698175906
transform 1 0 4928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698175906
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_37
timestamp 1698175906
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_45
timestamp 1698175906
transform 1 0 6384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_49
timestamp 1698175906
transform 1 0 6832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_58
timestamp 1698175906
transform 1 0 7840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_62
timestamp 1698175906
transform 1 0 8288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_64
timestamp 1698175906
transform 1 0 8512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_102
timestamp 1698175906
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698175906
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_115
timestamp 1698175906
transform 1 0 14224 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_131
timestamp 1698175906
transform 1 0 16016 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_139
timestamp 1698175906
transform 1 0 16912 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_143
timestamp 1698175906
transform 1 0 17360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_152
timestamp 1698175906
transform 1 0 18368 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_168
timestamp 1698175906
transform 1 0 20160 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_172
timestamp 1698175906
transform 1 0 20608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698175906
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_185
timestamp 1698175906
transform 1 0 22064 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_191
timestamp 1698175906
transform 1 0 22736 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_193
timestamp 1698175906
transform 1 0 22960 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_196
timestamp 1698175906
transform 1 0 23296 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_202
timestamp 1698175906
transform 1 0 23968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_211
timestamp 1698175906
transform 1 0 24976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_243
timestamp 1698175906
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698175906
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_295
timestamp 1698175906
transform 1 0 34384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_297
timestamp 1698175906
transform 1 0 34608 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_300
timestamp 1698175906
transform 1 0 34944 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_308
timestamp 1698175906
transform 1 0 35840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_312
timestamp 1698175906
transform 1 0 36288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698175906
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_317
timestamp 1698175906
transform 1 0 36848 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_333
timestamp 1698175906
transform 1 0 38640 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_341
timestamp 1698175906
transform 1 0 39536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_345
timestamp 1698175906
transform 1 0 39984 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_356
timestamp 1698175906
transform 1 0 41216 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_372
timestamp 1698175906
transform 1 0 43008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_380
timestamp 1698175906
transform 1 0 43904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_384
timestamp 1698175906
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698175906
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698175906
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_457
timestamp 1698175906
transform 1 0 52528 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_489
timestamp 1698175906
transform 1 0 56112 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_505
timestamp 1698175906
transform 1 0 57904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1698175906
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_6
timestamp 1698175906
transform 1 0 2016 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_16
timestamp 1698175906
transform 1 0 3136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_105
timestamp 1698175906
transform 1 0 13104 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_109
timestamp 1698175906
transform 1 0 13552 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_119
timestamp 1698175906
transform 1 0 14672 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_135
timestamp 1698175906
transform 1 0 16464 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698175906
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_189
timestamp 1698175906
transform 1 0 22512 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_193
timestamp 1698175906
transform 1 0 22960 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_204
timestamp 1698175906
transform 1 0 24192 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_212
timestamp 1698175906
transform 1 0 25088 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_267
timestamp 1698175906
transform 1 0 31248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_269
timestamp 1698175906
transform 1 0 31472 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_276
timestamp 1698175906
transform 1 0 32256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_288
timestamp 1698175906
transform 1 0 33600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_318
timestamp 1698175906
transform 1 0 36960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_324
timestamp 1698175906
transform 1 0 37632 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_344
timestamp 1698175906
transform 1 0 39872 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698175906
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698175906
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_362
timestamp 1698175906
transform 1 0 41888 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_394
timestamp 1698175906
transform 1 0 45472 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_410
timestamp 1698175906
transform 1 0 47264 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_418
timestamp 1698175906
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698175906
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698175906
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698175906
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698175906
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698175906
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698175906
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_51
timestamp 1698175906
transform 1 0 7056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_67
timestamp 1698175906
transform 1 0 8848 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_71
timestamp 1698175906
transform 1 0 9296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_73
timestamp 1698175906
transform 1 0 9520 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698175906
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698175906
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_111
timestamp 1698175906
transform 1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_113
timestamp 1698175906
transform 1 0 14000 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_130
timestamp 1698175906
transform 1 0 15904 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_177
timestamp 1698175906
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_181
timestamp 1698175906
transform 1 0 21616 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_189
timestamp 1698175906
transform 1 0 22512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_200
timestamp 1698175906
transform 1 0 23744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_204
timestamp 1698175906
transform 1 0 24192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_207
timestamp 1698175906
transform 1 0 24528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_231
timestamp 1698175906
transform 1 0 27216 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_242
timestamp 1698175906
transform 1 0 28448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698175906
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_257
timestamp 1698175906
transform 1 0 30128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_259
timestamp 1698175906
transform 1 0 30352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_302
timestamp 1698175906
transform 1 0 35168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_306
timestamp 1698175906
transform 1 0 35616 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698175906
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_317
timestamp 1698175906
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_348
timestamp 1698175906
transform 1 0 40320 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_358
timestamp 1698175906
transform 1 0 41440 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_374
timestamp 1698175906
transform 1 0 43232 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_382
timestamp 1698175906
transform 1 0 44128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698175906
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_387
timestamp 1698175906
transform 1 0 44688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698175906
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_457
timestamp 1698175906
transform 1 0 52528 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_489
timestamp 1698175906
transform 1 0 56112 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_505
timestamp 1698175906
transform 1 0 57904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2
timestamp 1698175906
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_6
timestamp 1698175906
transform 1 0 2016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_8
timestamp 1698175906
transform 1 0 2240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_19
timestamp 1698175906
transform 1 0 3472 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_28
timestamp 1698175906
transform 1 0 4480 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_64
timestamp 1698175906
transform 1 0 8512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698175906
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_72
timestamp 1698175906
transform 1 0 9408 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_99
timestamp 1698175906
transform 1 0 12432 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_107
timestamp 1698175906
transform 1 0 13328 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_117
timestamp 1698175906
transform 1 0 14448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_133
timestamp 1698175906
transform 1 0 16240 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_137
timestamp 1698175906
transform 1 0 16688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_139
timestamp 1698175906
transform 1 0 16912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_142
timestamp 1698175906
transform 1 0 17248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_150
timestamp 1698175906
transform 1 0 18144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_152
timestamp 1698175906
transform 1 0 18368 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_198
timestamp 1698175906
transform 1 0 23520 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_206
timestamp 1698175906
transform 1 0 24416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698175906
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_216
timestamp 1698175906
transform 1 0 25536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_257
timestamp 1698175906
transform 1 0 30128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_261
timestamp 1698175906
transform 1 0 30576 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_277
timestamp 1698175906
transform 1 0 32368 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698175906
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_284
timestamp 1698175906
transform 1 0 33152 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_343
timestamp 1698175906
transform 1 0 39760 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_347
timestamp 1698175906
transform 1 0 40208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698175906
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_352
timestamp 1698175906
transform 1 0 40768 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_356
timestamp 1698175906
transform 1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_387
timestamp 1698175906
transform 1 0 44688 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698175906
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698175906
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698175906
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698175906
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698175906
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_8
timestamp 1698175906
transform 1 0 2240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_12
timestamp 1698175906
transform 1 0 2688 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_20
timestamp 1698175906
transform 1 0 3584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_30
timestamp 1698175906
transform 1 0 4704 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698175906
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_37
timestamp 1698175906
transform 1 0 5488 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_67
timestamp 1698175906
transform 1 0 8848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_69
timestamp 1698175906
transform 1 0 9072 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_78
timestamp 1698175906
transform 1 0 10080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_107
timestamp 1698175906
transform 1 0 13328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_119
timestamp 1698175906
transform 1 0 14672 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_127
timestamp 1698175906
transform 1 0 15568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_139
timestamp 1698175906
transform 1 0 16912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_143
timestamp 1698175906
transform 1 0 17360 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_147
timestamp 1698175906
transform 1 0 17808 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_169
timestamp 1698175906
transform 1 0 20272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_173
timestamp 1698175906
transform 1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698175906
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_190
timestamp 1698175906
transform 1 0 22624 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_194
timestamp 1698175906
transform 1 0 23072 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_301
timestamp 1698175906
transform 1 0 35056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_309
timestamp 1698175906
transform 1 0 35952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1698175906
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_317
timestamp 1698175906
transform 1 0 36848 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_335
timestamp 1698175906
transform 1 0 38864 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_351
timestamp 1698175906
transform 1 0 40656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_353
timestamp 1698175906
transform 1 0 40880 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_364
timestamp 1698175906
transform 1 0 42112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_380
timestamp 1698175906
transform 1 0 43904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698175906
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_387
timestamp 1698175906
transform 1 0 44688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698175906
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_457
timestamp 1698175906
transform 1 0 52528 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_489
timestamp 1698175906
transform 1 0 56112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_505
timestamp 1698175906
transform 1 0 57904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_8
timestamp 1698175906
transform 1 0 2240 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_12
timestamp 1698175906
transform 1 0 2688 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_26
timestamp 1698175906
transform 1 0 4256 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_72
timestamp 1698175906
transform 1 0 9408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_126
timestamp 1698175906
transform 1 0 15456 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_130
timestamp 1698175906
transform 1 0 15904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_134
timestamp 1698175906
transform 1 0 16352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_138
timestamp 1698175906
transform 1 0 16800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_142
timestamp 1698175906
transform 1 0 17248 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_158
timestamp 1698175906
transform 1 0 19040 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_166
timestamp 1698175906
transform 1 0 19936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_170
timestamp 1698175906
transform 1 0 20384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_197
timestamp 1698175906
transform 1 0 23408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_201
timestamp 1698175906
transform 1 0 23856 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_203
timestamp 1698175906
transform 1 0 24080 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_206
timestamp 1698175906
transform 1 0 24416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_262
timestamp 1698175906
transform 1 0 30688 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_290
timestamp 1698175906
transform 1 0 33824 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_294
timestamp 1698175906
transform 1 0 34272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_324
timestamp 1698175906
transform 1 0 37632 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_328
timestamp 1698175906
transform 1 0 38080 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_342
timestamp 1698175906
transform 1 0 39648 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_346
timestamp 1698175906
transform 1 0 40096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_360
timestamp 1698175906
transform 1 0 41664 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_392
timestamp 1698175906
transform 1 0 45248 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_408
timestamp 1698175906
transform 1 0 47040 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698175906
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_422
timestamp 1698175906
transform 1 0 48608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698175906
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698175906
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698175906
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2
timestamp 1698175906
transform 1 0 1568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_30
timestamp 1698175906
transform 1 0 4704 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698175906
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_37
timestamp 1698175906
transform 1 0 5488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_41
timestamp 1698175906
transform 1 0 5936 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_50
timestamp 1698175906
transform 1 0 6944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_133
timestamp 1698175906
transform 1 0 16240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_137
timestamp 1698175906
transform 1 0 16688 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_139
timestamp 1698175906
transform 1 0 16912 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_145
timestamp 1698175906
transform 1 0 17584 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_157
timestamp 1698175906
transform 1 0 18928 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698175906
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_177
timestamp 1698175906
transform 1 0 21168 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_209
timestamp 1698175906
transform 1 0 24752 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_279
timestamp 1698175906
transform 1 0 32592 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_291
timestamp 1698175906
transform 1 0 33936 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_295
timestamp 1698175906
transform 1 0 34384 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_304
timestamp 1698175906
transform 1 0 35392 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_308
timestamp 1698175906
transform 1 0 35840 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_312
timestamp 1698175906
transform 1 0 36288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698175906
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_317
timestamp 1698175906
transform 1 0 36848 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_325
timestamp 1698175906
transform 1 0 37744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_327
timestamp 1698175906
transform 1 0 37968 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_373
timestamp 1698175906
transform 1 0 43120 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_381
timestamp 1698175906
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_387
timestamp 1698175906
transform 1 0 44688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698175906
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_457
timestamp 1698175906
transform 1 0 52528 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_489
timestamp 1698175906
transform 1 0 56112 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_505
timestamp 1698175906
transform 1 0 57904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_2
timestamp 1698175906
transform 1 0 1568 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_26
timestamp 1698175906
transform 1 0 4256 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_34
timestamp 1698175906
transform 1 0 5152 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_38
timestamp 1698175906
transform 1 0 5600 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_40
timestamp 1698175906
transform 1 0 5824 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_54
timestamp 1698175906
transform 1 0 7392 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_72
timestamp 1698175906
transform 1 0 9408 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_97
timestamp 1698175906
transform 1 0 12208 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_105
timestamp 1698175906
transform 1 0 13104 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_118
timestamp 1698175906
transform 1 0 14560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_130
timestamp 1698175906
transform 1 0 15904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_132
timestamp 1698175906
transform 1 0 16128 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_135
timestamp 1698175906
transform 1 0 16464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_139
timestamp 1698175906
transform 1 0 16912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_169
timestamp 1698175906
transform 1 0 20272 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_173
timestamp 1698175906
transform 1 0 20720 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_177
timestamp 1698175906
transform 1 0 21168 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_185
timestamp 1698175906
transform 1 0 22064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_187
timestamp 1698175906
transform 1 0 22288 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_205
timestamp 1698175906
transform 1 0 24304 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698175906
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_212
timestamp 1698175906
transform 1 0 25088 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_220
timestamp 1698175906
transform 1 0 25984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_222
timestamp 1698175906
transform 1 0 26208 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_273
timestamp 1698175906
transform 1 0 31920 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_277
timestamp 1698175906
transform 1 0 32368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698175906
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_282
timestamp 1698175906
transform 1 0 32928 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_339
timestamp 1698175906
transform 1 0 39312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_341
timestamp 1698175906
transform 1 0 39536 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_344
timestamp 1698175906
transform 1 0 39872 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_348
timestamp 1698175906
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_352
timestamp 1698175906
transform 1 0 40768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698175906
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698175906
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698175906
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698175906
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698175906
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_8
timestamp 1698175906
transform 1 0 2240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_12
timestamp 1698175906
transform 1 0 2688 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_28
timestamp 1698175906
transform 1 0 4480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698175906
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698175906
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_37
timestamp 1698175906
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_53
timestamp 1698175906
transform 1 0 7280 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_69
timestamp 1698175906
transform 1 0 9072 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_81
timestamp 1698175906
transform 1 0 10416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_85
timestamp 1698175906
transform 1 0 10864 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_92
timestamp 1698175906
transform 1 0 11648 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_96
timestamp 1698175906
transform 1 0 12096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_98
timestamp 1698175906
transform 1 0 12320 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698175906
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_107
timestamp 1698175906
transform 1 0 13328 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_118
timestamp 1698175906
transform 1 0 14560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_137
timestamp 1698175906
transform 1 0 16688 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_141
timestamp 1698175906
transform 1 0 17136 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_154
timestamp 1698175906
transform 1 0 18592 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_173
timestamp 1698175906
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_177
timestamp 1698175906
transform 1 0 21168 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_196
timestamp 1698175906
transform 1 0 23296 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_204
timestamp 1698175906
transform 1 0 24192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_242
timestamp 1698175906
transform 1 0 28448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698175906
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_247
timestamp 1698175906
transform 1 0 29008 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_288
timestamp 1698175906
transform 1 0 33600 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_308
timestamp 1698175906
transform 1 0 35840 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_312
timestamp 1698175906
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698175906
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_317
timestamp 1698175906
transform 1 0 36848 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_325
timestamp 1698175906
transform 1 0 37744 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_329
timestamp 1698175906
transform 1 0 38192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_333
timestamp 1698175906
transform 1 0 38640 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_365
timestamp 1698175906
transform 1 0 42224 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698175906
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698175906
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698175906
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_457
timestamp 1698175906
transform 1 0 52528 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_489
timestamp 1698175906
transform 1 0 56112 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_505
timestamp 1698175906
transform 1 0 57904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_31
timestamp 1698175906
transform 1 0 4816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_35
timestamp 1698175906
transform 1 0 5264 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_39
timestamp 1698175906
transform 1 0 5712 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_72
timestamp 1698175906
transform 1 0 9408 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_84
timestamp 1698175906
transform 1 0 10752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_86
timestamp 1698175906
transform 1 0 10976 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_99
timestamp 1698175906
transform 1 0 12432 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_107
timestamp 1698175906
transform 1 0 13328 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_115
timestamp 1698175906
transform 1 0 14224 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_119
timestamp 1698175906
transform 1 0 14672 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_122
timestamp 1698175906
transform 1 0 15008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_126
timestamp 1698175906
transform 1 0 15456 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_134
timestamp 1698175906
transform 1 0 16352 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_138
timestamp 1698175906
transform 1 0 16800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_142
timestamp 1698175906
transform 1 0 17248 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_174
timestamp 1698175906
transform 1 0 20832 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_190
timestamp 1698175906
transform 1 0 22624 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698175906
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_216
timestamp 1698175906
transform 1 0 25536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_220
timestamp 1698175906
transform 1 0 25984 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_228
timestamp 1698175906
transform 1 0 26880 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_232
timestamp 1698175906
transform 1 0 27328 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_237
timestamp 1698175906
transform 1 0 27888 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_245
timestamp 1698175906
transform 1 0 28784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_247
timestamp 1698175906
transform 1 0 29008 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_277
timestamp 1698175906
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698175906
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_282
timestamp 1698175906
transform 1 0 32928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_286
timestamp 1698175906
transform 1 0 33376 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_323
timestamp 1698175906
transform 1 0 37520 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_327
timestamp 1698175906
transform 1 0 37968 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_343
timestamp 1698175906
transform 1 0 39760 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_347
timestamp 1698175906
transform 1 0 40208 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698175906
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_352
timestamp 1698175906
transform 1 0 40768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698175906
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698175906
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698175906
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698175906
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698175906
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_31
timestamp 1698175906
transform 1 0 4816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_37
timestamp 1698175906
transform 1 0 5488 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_45
timestamp 1698175906
transform 1 0 6384 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_49
timestamp 1698175906
transform 1 0 6832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_58
timestamp 1698175906
transform 1 0 7840 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_90
timestamp 1698175906
transform 1 0 11424 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_92
timestamp 1698175906
transform 1 0 11648 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_95
timestamp 1698175906
transform 1 0 11984 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698175906
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_107
timestamp 1698175906
transform 1 0 13328 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_123
timestamp 1698175906
transform 1 0 15120 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_127
timestamp 1698175906
transform 1 0 15568 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_133
timestamp 1698175906
transform 1 0 16240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_137
timestamp 1698175906
transform 1 0 16688 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_141
timestamp 1698175906
transform 1 0 17136 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_148
timestamp 1698175906
transform 1 0 17920 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_157
timestamp 1698175906
transform 1 0 18928 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_173
timestamp 1698175906
transform 1 0 20720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_220
timestamp 1698175906
transform 1 0 25984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_230
timestamp 1698175906
transform 1 0 27104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_234
timestamp 1698175906
transform 1 0 27552 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_242
timestamp 1698175906
transform 1 0 28448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698175906
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_247
timestamp 1698175906
transform 1 0 29008 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_255
timestamp 1698175906
transform 1 0 29904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_263
timestamp 1698175906
transform 1 0 30800 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_271
timestamp 1698175906
transform 1 0 31696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_275
timestamp 1698175906
transform 1 0 32144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_279
timestamp 1698175906
transform 1 0 32592 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_295
timestamp 1698175906
transform 1 0 34384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_305
timestamp 1698175906
transform 1 0 35504 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_317
timestamp 1698175906
transform 1 0 36848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_348
timestamp 1698175906
transform 1 0 40320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_352
timestamp 1698175906
transform 1 0 40768 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698175906
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698175906
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698175906
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_457
timestamp 1698175906
transform 1 0 52528 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_489
timestamp 1698175906
transform 1 0 56112 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_505
timestamp 1698175906
transform 1 0 57904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_8
timestamp 1698175906
transform 1 0 2240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_12
timestamp 1698175906
transform 1 0 2688 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_20
timestamp 1698175906
transform 1 0 3584 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_24
timestamp 1698175906
transform 1 0 4032 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_54
timestamp 1698175906
transform 1 0 7392 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_58
timestamp 1698175906
transform 1 0 7840 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698175906
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_72
timestamp 1698175906
transform 1 0 9408 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_80
timestamp 1698175906
transform 1 0 10304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_92
timestamp 1698175906
transform 1 0 11648 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_96
timestamp 1698175906
transform 1 0 12096 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_133
timestamp 1698175906
transform 1 0 16240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_192
timestamp 1698175906
transform 1 0 22848 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_196
timestamp 1698175906
transform 1 0 23296 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_204
timestamp 1698175906
transform 1 0 24192 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_208
timestamp 1698175906
transform 1 0 24640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_212
timestamp 1698175906
transform 1 0 25088 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_242
timestamp 1698175906
transform 1 0 28448 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_274
timestamp 1698175906
transform 1 0 32032 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_278
timestamp 1698175906
transform 1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_282
timestamp 1698175906
transform 1 0 32928 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_298
timestamp 1698175906
transform 1 0 34720 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_306
timestamp 1698175906
transform 1 0 35616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_310
timestamp 1698175906
transform 1 0 36064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_312
timestamp 1698175906
transform 1 0 36288 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_315
timestamp 1698175906
transform 1 0 36624 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_331
timestamp 1698175906
transform 1 0 38416 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_352
timestamp 1698175906
transform 1 0 40768 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_369
timestamp 1698175906
transform 1 0 42672 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_401
timestamp 1698175906
transform 1 0 46256 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_417
timestamp 1698175906
transform 1 0 48048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_419
timestamp 1698175906
transform 1 0 48272 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698175906
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698175906
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698175906
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698175906
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698175906
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698175906
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_37
timestamp 1698175906
transform 1 0 5488 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_53
timestamp 1698175906
transform 1 0 7280 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_61
timestamp 1698175906
transform 1 0 8176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_65
timestamp 1698175906
transform 1 0 8624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_67
timestamp 1698175906
transform 1 0 8848 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_70
timestamp 1698175906
transform 1 0 9184 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_74
timestamp 1698175906
transform 1 0 9632 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_96
timestamp 1698175906
transform 1 0 12096 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_100
timestamp 1698175906
transform 1 0 12544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_104
timestamp 1698175906
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_107
timestamp 1698175906
transform 1 0 13328 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_115
timestamp 1698175906
transform 1 0 14224 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_133
timestamp 1698175906
transform 1 0 16240 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_141
timestamp 1698175906
transform 1 0 17136 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_145
timestamp 1698175906
transform 1 0 17584 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_177
timestamp 1698175906
transform 1 0 21168 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_231
timestamp 1698175906
transform 1 0 27216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_235
timestamp 1698175906
transform 1 0 27664 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_243
timestamp 1698175906
transform 1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_247
timestamp 1698175906
transform 1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_278
timestamp 1698175906
transform 1 0 32480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_282
timestamp 1698175906
transform 1 0 32928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1698175906
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_323
timestamp 1698175906
transform 1 0 37520 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_327
timestamp 1698175906
transform 1 0 37968 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_354
timestamp 1698175906
transform 1 0 40992 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_358
timestamp 1698175906
transform 1 0 41440 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_362
timestamp 1698175906
transform 1 0 41888 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_378
timestamp 1698175906
transform 1 0 43680 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_382
timestamp 1698175906
transform 1 0 44128 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_384
timestamp 1698175906
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698175906
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698175906
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698175906
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698175906
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698175906
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_8
timestamp 1698175906
transform 1 0 2240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_12
timestamp 1698175906
transform 1 0 2688 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_28
timestamp 1698175906
transform 1 0 4480 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_36
timestamp 1698175906
transform 1 0 5376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_38
timestamp 1698175906
transform 1 0 5600 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_68
timestamp 1698175906
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_72
timestamp 1698175906
transform 1 0 9408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_74
timestamp 1698175906
transform 1 0 9632 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_91
timestamp 1698175906
transform 1 0 11536 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_93
timestamp 1698175906
transform 1 0 11760 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_100
timestamp 1698175906
transform 1 0 12544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_104
timestamp 1698175906
transform 1 0 12992 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_120
timestamp 1698175906
transform 1 0 14784 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_124
timestamp 1698175906
transform 1 0 15232 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_127
timestamp 1698175906
transform 1 0 15568 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_135
timestamp 1698175906
transform 1 0 16464 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698175906
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_142
timestamp 1698175906
transform 1 0 17248 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_146
timestamp 1698175906
transform 1 0 17696 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_156
timestamp 1698175906
transform 1 0 18816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_160
timestamp 1698175906
transform 1 0 19264 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_176
timestamp 1698175906
transform 1 0 21056 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_184
timestamp 1698175906
transform 1 0 21952 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_186
timestamp 1698175906
transform 1 0 22176 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_195
timestamp 1698175906
transform 1 0 23184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_199
timestamp 1698175906
transform 1 0 23632 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_207
timestamp 1698175906
transform 1 0 24528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_209
timestamp 1698175906
transform 1 0 24752 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698175906
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_214
timestamp 1698175906
transform 1 0 25312 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_223
timestamp 1698175906
transform 1 0 26320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_231
timestamp 1698175906
transform 1 0 27216 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_235
timestamp 1698175906
transform 1 0 27664 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_243
timestamp 1698175906
transform 1 0 28560 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_247
timestamp 1698175906
transform 1 0 29008 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_264
timestamp 1698175906
transform 1 0 30912 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_268
timestamp 1698175906
transform 1 0 31360 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_270
timestamp 1698175906
transform 1 0 31584 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_277
timestamp 1698175906
transform 1 0 32368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_279
timestamp 1698175906
transform 1 0 32592 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_292
timestamp 1698175906
transform 1 0 34048 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_308
timestamp 1698175906
transform 1 0 35840 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_321
timestamp 1698175906
transform 1 0 37296 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_337
timestamp 1698175906
transform 1 0 39088 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_345
timestamp 1698175906
transform 1 0 39984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_347
timestamp 1698175906
transform 1 0 40208 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_391
timestamp 1698175906
transform 1 0 45136 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_407
timestamp 1698175906
transform 1 0 46928 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_415
timestamp 1698175906
transform 1 0 47824 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_419
timestamp 1698175906
transform 1 0 48272 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698175906
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698175906
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698175906
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698175906
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698175906
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698175906
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_37
timestamp 1698175906
transform 1 0 5488 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_69
timestamp 1698175906
transform 1 0 9072 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_77
timestamp 1698175906
transform 1 0 9968 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_83
timestamp 1698175906
transform 1 0 10640 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_93
timestamp 1698175906
transform 1 0 11760 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698175906
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_107
timestamp 1698175906
transform 1 0 13328 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_123
timestamp 1698175906
transform 1 0 15120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_127
timestamp 1698175906
transform 1 0 15568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_129
timestamp 1698175906
transform 1 0 15792 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_138
timestamp 1698175906
transform 1 0 16800 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_146
timestamp 1698175906
transform 1 0 17696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_152
timestamp 1698175906
transform 1 0 18368 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_168
timestamp 1698175906
transform 1 0 20160 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_172
timestamp 1698175906
transform 1 0 20608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698175906
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_177
timestamp 1698175906
transform 1 0 21168 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_181
timestamp 1698175906
transform 1 0 21616 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_183
timestamp 1698175906
transform 1 0 21840 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_194
timestamp 1698175906
transform 1 0 23072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_196
timestamp 1698175906
transform 1 0 23296 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_205
timestamp 1698175906
transform 1 0 24304 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_214
timestamp 1698175906
transform 1 0 25312 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_218
timestamp 1698175906
transform 1 0 25760 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_220
timestamp 1698175906
transform 1 0 25984 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_229
timestamp 1698175906
transform 1 0 26992 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_247
timestamp 1698175906
transform 1 0 29008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_251
timestamp 1698175906
transform 1 0 29456 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_267
timestamp 1698175906
transform 1 0 31248 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_275
timestamp 1698175906
transform 1 0 32144 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_287
timestamp 1698175906
transform 1 0 33488 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_303
timestamp 1698175906
transform 1 0 35280 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698175906
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_317
timestamp 1698175906
transform 1 0 36848 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_321
timestamp 1698175906
transform 1 0 37296 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_323
timestamp 1698175906
transform 1 0 37520 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_332
timestamp 1698175906
transform 1 0 38528 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_334
timestamp 1698175906
transform 1 0 38752 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_337
timestamp 1698175906
transform 1 0 39088 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_345
timestamp 1698175906
transform 1 0 39984 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_349
timestamp 1698175906
transform 1 0 40432 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_351
timestamp 1698175906
transform 1 0 40656 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_358
timestamp 1698175906
transform 1 0 41440 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_368
timestamp 1698175906
transform 1 0 42560 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1698175906
transform 1 0 44352 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698175906
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698175906
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698175906
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698175906
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698175906
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_8
timestamp 1698175906
transform 1 0 2240 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_12
timestamp 1698175906
transform 1 0 2688 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_44
timestamp 1698175906
transform 1 0 6272 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_60
timestamp 1698175906
transform 1 0 8064 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_68
timestamp 1698175906
transform 1 0 8960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_72
timestamp 1698175906
transform 1 0 9408 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_88
timestamp 1698175906
transform 1 0 11200 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_96
timestamp 1698175906
transform 1 0 12096 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_113
timestamp 1698175906
transform 1 0 14000 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_125
timestamp 1698175906
transform 1 0 15344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_135
timestamp 1698175906
transform 1 0 16464 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_139
timestamp 1698175906
transform 1 0 16912 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_158
timestamp 1698175906
transform 1 0 19040 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_203
timestamp 1698175906
transform 1 0 24080 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_207
timestamp 1698175906
transform 1 0 24528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698175906
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_241
timestamp 1698175906
transform 1 0 28336 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_263
timestamp 1698175906
transform 1 0 30800 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_267
timestamp 1698175906
transform 1 0 31248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_269
timestamp 1698175906
transform 1 0 31472 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_276
timestamp 1698175906
transform 1 0 32256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_282
timestamp 1698175906
transform 1 0 32928 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_293
timestamp 1698175906
transform 1 0 34160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_295
timestamp 1698175906
transform 1 0 34384 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_302
timestamp 1698175906
transform 1 0 35168 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_306
timestamp 1698175906
transform 1 0 35616 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_308
timestamp 1698175906
transform 1 0 35840 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_315
timestamp 1698175906
transform 1 0 36624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_319
timestamp 1698175906
transform 1 0 37072 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_327
timestamp 1698175906
transform 1 0 37968 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_343
timestamp 1698175906
transform 1 0 39760 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_347
timestamp 1698175906
transform 1 0 40208 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_362
timestamp 1698175906
transform 1 0 41888 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_394
timestamp 1698175906
transform 1 0 45472 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_410
timestamp 1698175906
transform 1 0 47264 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_418
timestamp 1698175906
transform 1 0 48160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_422
timestamp 1698175906
transform 1 0 48608 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_454
timestamp 1698175906
transform 1 0 52192 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_470
timestamp 1698175906
transform 1 0 53984 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_478
timestamp 1698175906
transform 1 0 54880 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_480
timestamp 1698175906
transform 1 0 55104 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_483
timestamp 1698175906
transform 1 0 55440 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_487
timestamp 1698175906
transform 1 0 55888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_489
timestamp 1698175906
transform 1 0 56112 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698175906
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698175906
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2
timestamp 1698175906
transform 1 0 1568 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_8
timestamp 1698175906
transform 1 0 2240 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_24
timestamp 1698175906
transform 1 0 4032 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698175906
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698175906
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_37
timestamp 1698175906
transform 1 0 5488 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_69
timestamp 1698175906
transform 1 0 9072 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_85
timestamp 1698175906
transform 1 0 10864 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_89
timestamp 1698175906
transform 1 0 11312 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_91
timestamp 1698175906
transform 1 0 11536 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_96
timestamp 1698175906
transform 1 0 12096 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_104
timestamp 1698175906
transform 1 0 12992 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_136
timestamp 1698175906
transform 1 0 16576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_140
timestamp 1698175906
transform 1 0 17024 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_173
timestamp 1698175906
transform 1 0 20720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_177
timestamp 1698175906
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_181
timestamp 1698175906
transform 1 0 21616 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_189
timestamp 1698175906
transform 1 0 22512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_195
timestamp 1698175906
transform 1 0 23184 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_211
timestamp 1698175906
transform 1 0 24976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_217
timestamp 1698175906
transform 1 0 25648 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_237
timestamp 1698175906
transform 1 0 27888 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_282
timestamp 1698175906
transform 1 0 32928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_323
timestamp 1698175906
transform 1 0 37520 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_339
timestamp 1698175906
transform 1 0 39312 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_343
timestamp 1698175906
transform 1 0 39760 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_375
timestamp 1698175906
transform 1 0 43344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_379
timestamp 1698175906
transform 1 0 43792 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_383
timestamp 1698175906
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_387
timestamp 1698175906
transform 1 0 44688 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_391
timestamp 1698175906
transform 1 0 45136 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_421
timestamp 1698175906
transform 1 0 48496 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_437
timestamp 1698175906
transform 1 0 50288 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_441
timestamp 1698175906
transform 1 0 50736 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_444
timestamp 1698175906
transform 1 0 51072 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_452
timestamp 1698175906
transform 1 0 51968 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_14
timestamp 1698175906
transform 1 0 2912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1698175906
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_26
timestamp 1698175906
transform 1 0 4256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_30
timestamp 1698175906
transform 1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_42
timestamp 1698175906
transform 1 0 6048 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_50
timestamp 1698175906
transform 1 0 6944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_52
timestamp 1698175906
transform 1 0 7168 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_61
timestamp 1698175906
transform 1 0 8176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_65
timestamp 1698175906
transform 1 0 8624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_67
timestamp 1698175906
transform 1 0 8848 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_70
timestamp 1698175906
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_72
timestamp 1698175906
transform 1 0 9408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_81
timestamp 1698175906
transform 1 0 10416 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_89
timestamp 1698175906
transform 1 0 11312 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_101
timestamp 1698175906
transform 1 0 12656 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_104
timestamp 1698175906
transform 1 0 12992 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_112
timestamp 1698175906
transform 1 0 13888 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_121
timestamp 1698175906
transform 1 0 14896 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_129
timestamp 1698175906
transform 1 0 15792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_133
timestamp 1698175906
transform 1 0 16240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_144
timestamp 1698175906
transform 1 0 17472 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_152
timestamp 1698175906
transform 1 0 18368 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_161
timestamp 1698175906
transform 1 0 19376 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_165
timestamp 1698175906
transform 1 0 19824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_167
timestamp 1698175906
transform 1 0 20048 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_172
timestamp 1698175906
transform 1 0 20608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_174
timestamp 1698175906
transform 1 0 20832 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_181
timestamp 1698175906
transform 1 0 21616 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_189
timestamp 1698175906
transform 1 0 22512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_201
timestamp 1698175906
transform 1 0 23856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_203
timestamp 1698175906
transform 1 0 24080 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698175906
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_210
timestamp 1698175906
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_212
timestamp 1698175906
transform 1 0 25088 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_221
timestamp 1698175906
transform 1 0 26096 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_229
timestamp 1698175906
transform 1 0 26992 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_233
timestamp 1698175906
transform 1 0 27440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_235
timestamp 1698175906
transform 1 0 27664 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_246
timestamp 1698175906
transform 1 0 28896 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_250
timestamp 1698175906
transform 1 0 29344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_252
timestamp 1698175906
transform 1 0 29568 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_261
timestamp 1698175906
transform 1 0 30576 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_269
timestamp 1698175906
transform 1 0 31472 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_274
timestamp 1698175906
transform 1 0 32032 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_281
timestamp 1698175906
transform 1 0 32816 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_289
timestamp 1698175906
transform 1 0 33712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_301
timestamp 1698175906
transform 1 0 35056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_305
timestamp 1698175906
transform 1 0 35504 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_308
timestamp 1698175906
transform 1 0 35840 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_312
timestamp 1698175906
transform 1 0 36288 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_321
timestamp 1698175906
transform 1 0 37296 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_329
timestamp 1698175906
transform 1 0 38192 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_333
timestamp 1698175906
transform 1 0 38640 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_336
timestamp 1698175906
transform 1 0 38976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_402
timestamp 1698175906
transform 1 0 46368 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_406
timestamp 1698175906
transform 1 0 46816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_410
timestamp 1698175906
transform 1 0 47264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_412
timestamp 1698175906
transform 1 0 47488 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698175906
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_470
timestamp 1698175906
transform 1 0 53984 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_504
timestamp 1698175906
transform 1 0 57792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698175906
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698175906
transform 1 0 7504 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698175906
transform -1 0 23856 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698175906
transform -1 0 26096 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698175906
transform -1 0 28896 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698175906
transform -1 0 30576 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698175906
transform 1 0 32144 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698175906
transform 1 0 34384 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698175906
transform 1 0 36624 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698175906
transform -1 0 40320 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698175906
transform 1 0 16800 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input11
timestamp 1698175906
transform 1 0 18704 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698175906
transform 1 0 20944 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1698175906
transform 1 0 11984 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698175906
transform 1 0 9744 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698175906
transform 1 0 1568 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698175906
transform 1 0 1568 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698175906
transform 1 0 1568 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698175906
transform 1 0 1568 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698175906
transform 1 0 1568 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698175906
transform -1 0 2912 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698175906
transform 1 0 1568 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698175906
transform 1 0 1568 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698175906
transform 1 0 1568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698175906
transform 1 0 1568 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698175906
transform 1 0 1568 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input31
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input32
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698175906
transform 1 0 2240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input39
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input45
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698175906
transform -1 0 14896 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698175906
transform 1 0 5376 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698175906
transform 1 0 43456 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698175906
transform 1 0 45584 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698175906
transform 1 0 47824 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698175906
transform 1 0 51072 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698175906
transform 1 0 52528 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698175906
transform 1 0 54880 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698175906
transform 1 0 55440 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698175906
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698175906
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698175906
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698175906
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698175906
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698175906
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698175906
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698175906
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698175906
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698175906
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698175906
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698175906
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698175906
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698175906
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698175906
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698175906
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698175906
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698175906
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698175906
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698175906
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698175906
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698175906
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698175906
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698175906
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698175906
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698175906
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698175906
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698175906
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698175906
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698175906
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698175906
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698175906
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698175906
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698175906
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698175906
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698175906
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698175906
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698175906
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698175906
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698175906
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698175906
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698175906
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698175906
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698175906
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698175906
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698175906
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698175906
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698175906
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698175906
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698175906
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698175906
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698175906
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698175906
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698175906
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698175906
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698175906
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698175906
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698175906
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698175906
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698175906
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698175906
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698175906
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698175906
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698175906
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698175906
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698175906
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698175906
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698175906
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698175906
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698175906
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698175906
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698175906
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698175906
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698175906
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698175906
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698175906
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698175906
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698175906
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698175906
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698175906
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698175906
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698175906
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698175906
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698175906
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698175906
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698175906
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698175906
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698175906
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698175906
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698175906
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698175906
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698175906
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698175906
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698175906
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698175906
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698175906
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698175906
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698175906
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698175906
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698175906
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698175906
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698175906
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698175906
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698175906
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698175906
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698175906
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698175906
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698175906
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698175906
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698175906
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698175906
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698175906
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698175906
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698175906
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698175906
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698175906
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698175906
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698175906
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698175906
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698175906
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698175906
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698175906
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698175906
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698175906
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698175906
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698175906
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698175906
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698175906
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698175906
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698175906
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698175906
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698175906
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698175906
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698175906
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698175906
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698175906
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698175906
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698175906
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698175906
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698175906
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698175906
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698175906
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698175906
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698175906
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698175906
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698175906
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698175906
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698175906
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698175906
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698175906
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698175906
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698175906
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698175906
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698175906
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698175906
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698175906
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698175906
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698175906
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698175906
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698175906
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698175906
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698175906
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698175906
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698175906
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698175906
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698175906
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698175906
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698175906
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698175906
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698175906
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698175906
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698175906
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698175906
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698175906
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698175906
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698175906
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698175906
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698175906
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698175906
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698175906
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698175906
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698175906
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698175906
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698175906
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698175906
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698175906
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698175906
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698175906
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698175906
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698175906
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698175906
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698175906
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698175906
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698175906
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698175906
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698175906
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698175906
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698175906
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698175906
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698175906
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698175906
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698175906
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698175906
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698175906
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698175906
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698175906
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698175906
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698175906
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698175906
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698175906
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698175906
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698175906
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698175906
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698175906
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698175906
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698175906
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698175906
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698175906
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698175906
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698175906
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698175906
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698175906
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698175906
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698175906
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698175906
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698175906
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698175906
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698175906
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698175906
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698175906
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698175906
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698175906
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698175906
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698175906
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698175906
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698175906
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698175906
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698175906
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698175906
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698175906
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698175906
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698175906
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698175906
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698175906
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698175906
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698175906
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698175906
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698175906
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698175906
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698175906
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698175906
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698175906
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698175906
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698175906
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698175906
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698175906
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698175906
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698175906
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698175906
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698175906
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698175906
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698175906
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698175906
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698175906
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698175906
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698175906
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698175906
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698175906
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698175906
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698175906
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698175906
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698175906
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698175906
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698175906
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698175906
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698175906
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698175906
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698175906
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698175906
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698175906
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698175906
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698175906
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698175906
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698175906
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698175906
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698175906
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698175906
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698175906
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698175906
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698175906
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698175906
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698175906
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698175906
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698175906
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698175906
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698175906
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698175906
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698175906
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698175906
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698175906
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698175906
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698175906
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698175906
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698175906
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698175906
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698175906
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698175906
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698175906
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698175906
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698175906
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698175906
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698175906
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698175906
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698175906
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698175906
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698175906
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698175906
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698175906
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698175906
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698175906
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698175906
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698175906
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698175906
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698175906
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698175906
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698175906
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698175906
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698175906
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698175906
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698175906
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698175906
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698175906
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
<< labels >>
flabel metal2 s 7392 59200 7504 60000 0 FreeSans 448 90 0 0 WEb_raw
port 0 nsew signal input
flabel metal2 s 23072 59200 23184 60000 0 FreeSans 448 90 0 0 bus_in[0]
port 1 nsew signal input
flabel metal2 s 25312 59200 25424 60000 0 FreeSans 448 90 0 0 bus_in[1]
port 2 nsew signal input
flabel metal2 s 27552 59200 27664 60000 0 FreeSans 448 90 0 0 bus_in[2]
port 3 nsew signal input
flabel metal2 s 29792 59200 29904 60000 0 FreeSans 448 90 0 0 bus_in[3]
port 4 nsew signal input
flabel metal2 s 32032 59200 32144 60000 0 FreeSans 448 90 0 0 bus_in[4]
port 5 nsew signal input
flabel metal2 s 34272 59200 34384 60000 0 FreeSans 448 90 0 0 bus_in[5]
port 6 nsew signal input
flabel metal2 s 36512 59200 36624 60000 0 FreeSans 448 90 0 0 bus_in[6]
port 7 nsew signal input
flabel metal2 s 38752 59200 38864 60000 0 FreeSans 448 90 0 0 bus_in[7]
port 8 nsew signal input
flabel metal2 s 40992 59200 41104 60000 0 FreeSans 448 90 0 0 bus_out[0]
port 9 nsew signal tristate
flabel metal2 s 43232 59200 43344 60000 0 FreeSans 448 90 0 0 bus_out[1]
port 10 nsew signal tristate
flabel metal2 s 45472 59200 45584 60000 0 FreeSans 448 90 0 0 bus_out[2]
port 11 nsew signal tristate
flabel metal2 s 47712 59200 47824 60000 0 FreeSans 448 90 0 0 bus_out[3]
port 12 nsew signal tristate
flabel metal2 s 49952 59200 50064 60000 0 FreeSans 448 90 0 0 bus_out[4]
port 13 nsew signal tristate
flabel metal2 s 52192 59200 52304 60000 0 FreeSans 448 90 0 0 bus_out[5]
port 14 nsew signal tristate
flabel metal2 s 54432 59200 54544 60000 0 FreeSans 448 90 0 0 bus_out[6]
port 15 nsew signal tristate
flabel metal2 s 56672 59200 56784 60000 0 FreeSans 448 90 0 0 bus_out[7]
port 16 nsew signal tristate
flabel metal2 s 16352 59200 16464 60000 0 FreeSans 448 90 0 0 cs_port[0]
port 17 nsew signal input
flabel metal2 s 18592 59200 18704 60000 0 FreeSans 448 90 0 0 cs_port[1]
port 18 nsew signal input
flabel metal2 s 20832 59200 20944 60000 0 FreeSans 448 90 0 0 cs_port[2]
port 19 nsew signal input
flabel metal2 s 11872 59200 11984 60000 0 FreeSans 448 90 0 0 le_hi_act
port 20 nsew signal input
flabel metal2 s 9632 59200 9744 60000 0 FreeSans 448 90 0 0 le_lo_act
port 21 nsew signal input
flabel metal3 s 0 30688 800 30800 0 FreeSans 448 0 0 0 ram_end[0]
port 22 nsew signal input
flabel metal3 s 0 48608 800 48720 0 FreeSans 448 0 0 0 ram_end[10]
port 23 nsew signal input
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 ram_end[11]
port 24 nsew signal input
flabel metal3 s 0 52192 800 52304 0 FreeSans 448 0 0 0 ram_end[12]
port 25 nsew signal input
flabel metal3 s 0 53984 800 54096 0 FreeSans 448 0 0 0 ram_end[13]
port 26 nsew signal input
flabel metal3 s 0 55776 800 55888 0 FreeSans 448 0 0 0 ram_end[14]
port 27 nsew signal input
flabel metal3 s 0 57568 800 57680 0 FreeSans 448 0 0 0 ram_end[15]
port 28 nsew signal input
flabel metal3 s 0 32480 800 32592 0 FreeSans 448 0 0 0 ram_end[1]
port 29 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 ram_end[2]
port 30 nsew signal input
flabel metal3 s 0 36064 800 36176 0 FreeSans 448 0 0 0 ram_end[3]
port 31 nsew signal input
flabel metal3 s 0 37856 800 37968 0 FreeSans 448 0 0 0 ram_end[4]
port 32 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 ram_end[5]
port 33 nsew signal input
flabel metal3 s 0 41440 800 41552 0 FreeSans 448 0 0 0 ram_end[6]
port 34 nsew signal input
flabel metal3 s 0 43232 800 43344 0 FreeSans 448 0 0 0 ram_end[7]
port 35 nsew signal input
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 ram_end[8]
port 36 nsew signal input
flabel metal3 s 0 46816 800 46928 0 FreeSans 448 0 0 0 ram_end[9]
port 37 nsew signal input
flabel metal3 s 0 2016 800 2128 0 FreeSans 448 0 0 0 ram_start[0]
port 38 nsew signal input
flabel metal3 s 0 19936 800 20048 0 FreeSans 448 0 0 0 ram_start[10]
port 39 nsew signal input
flabel metal3 s 0 21728 800 21840 0 FreeSans 448 0 0 0 ram_start[11]
port 40 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 ram_start[12]
port 41 nsew signal input
flabel metal3 s 0 25312 800 25424 0 FreeSans 448 0 0 0 ram_start[13]
port 42 nsew signal input
flabel metal3 s 0 27104 800 27216 0 FreeSans 448 0 0 0 ram_start[14]
port 43 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 ram_start[15]
port 44 nsew signal input
flabel metal3 s 0 3808 800 3920 0 FreeSans 448 0 0 0 ram_start[1]
port 45 nsew signal input
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 ram_start[2]
port 46 nsew signal input
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 ram_start[3]
port 47 nsew signal input
flabel metal3 s 0 9184 800 9296 0 FreeSans 448 0 0 0 ram_start[4]
port 48 nsew signal input
flabel metal3 s 0 10976 800 11088 0 FreeSans 448 0 0 0 ram_start[5]
port 49 nsew signal input
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 ram_start[6]
port 50 nsew signal input
flabel metal3 s 0 14560 800 14672 0 FreeSans 448 0 0 0 ram_start[7]
port 51 nsew signal input
flabel metal3 s 0 16352 800 16464 0 FreeSans 448 0 0 0 ram_start[8]
port 52 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 ram_start[9]
port 53 nsew signal input
flabel metal2 s 14112 59200 14224 60000 0 FreeSans 448 90 0 0 rom_enabled
port 54 nsew signal input
flabel metal2 s 5152 59200 5264 60000 0 FreeSans 448 90 0 0 rst
port 55 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 56 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 56 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 57 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 57 nsew ground bidirectional
flabel metal2 s 2912 59200 3024 60000 0 FreeSans 448 90 0 0 wb_clk_i
port 58 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 7448 57778 7448 57778 0 WEb_raw
rlabel metal3 7336 49896 7336 49896 0 _0000_
rlabel metal2 3864 51296 3864 51296 0 _0001_
rlabel metal3 9352 53032 9352 53032 0 _0002_
rlabel metal2 11928 51576 11928 51576 0 _0003_
rlabel metal2 37800 41608 37800 41608 0 _0004_
rlabel metal2 35784 40936 35784 40936 0 _0005_
rlabel metal3 37016 38920 37016 38920 0 _0006_
rlabel metal2 34664 43848 34664 43848 0 _0007_
rlabel metal2 22120 51128 22120 51128 0 _0008_
rlabel metal2 24808 53928 24808 53928 0 _0009_
rlabel metal3 22120 53704 22120 53704 0 _0010_
rlabel metal2 26488 50960 26488 50960 0 _0011_
rlabel metal2 41384 47096 41384 47096 0 _0012_
rlabel metal2 41720 41776 41720 41776 0 _0013_
rlabel metal2 39312 44408 39312 44408 0 _0014_
rlabel metal2 42392 45248 42392 45248 0 _0015_
rlabel metal2 29960 54936 29960 54936 0 _0016_
rlabel metal2 30128 52248 30128 52248 0 _0017_
rlabel metal2 34328 54936 34328 54936 0 _0018_
rlabel metal2 34104 52696 34104 52696 0 _0019_
rlabel metal2 38024 51128 38024 51128 0 _0020_
rlabel metal2 42840 53088 42840 53088 0 _0021_
rlabel metal3 41608 50456 41608 50456 0 _0022_
rlabel metal2 41048 54936 41048 54936 0 _0023_
rlabel metal2 14728 54936 14728 54936 0 _0024_
rlabel metal2 13944 51576 13944 51576 0 _0025_
rlabel metal2 17640 54768 17640 54768 0 _0026_
rlabel metal2 19992 52528 19992 52528 0 _0027_
rlabel metal2 31640 48440 31640 48440 0 _0028_
rlabel metal2 35560 49224 35560 49224 0 _0029_
rlabel metal3 35896 46760 35896 46760 0 _0030_
rlabel metal2 31416 49056 31416 49056 0 _0031_
rlabel metal2 27496 47992 27496 47992 0 _0032_
rlabel metal2 37240 52416 37240 52416 0 _0033_
rlabel metal3 40656 52024 40656 52024 0 _0034_
rlabel metal2 38696 52304 38696 52304 0 _0035_
rlabel metal2 37352 30184 37352 30184 0 _0036_
rlabel metal2 38248 37744 38248 37744 0 _0037_
rlabel metal2 33544 33488 33544 33488 0 _0038_
rlabel metal2 39256 33600 39256 33600 0 _0039_
rlabel metal2 35000 39200 35000 39200 0 _0040_
rlabel metal2 39704 31780 39704 31780 0 _0041_
rlabel metal3 32816 38808 32816 38808 0 _0042_
rlabel metal2 6664 47096 6664 47096 0 _0043_
rlabel metal3 5712 40488 5712 40488 0 _0044_
rlabel metal3 9520 47432 9520 47432 0 _0045_
rlabel metal2 11312 48216 11312 48216 0 _0046_
rlabel metal2 8344 47936 8344 47936 0 _0047_
rlabel metal2 12152 45808 12152 45808 0 _0048_
rlabel metal2 3976 47040 3976 47040 0 _0049_
rlabel metal3 6384 46760 6384 46760 0 _0050_
rlabel metal2 11704 48216 11704 48216 0 _0051_
rlabel metal2 14000 49000 14000 49000 0 _0052_
rlabel metal2 28168 44352 28168 44352 0 _0053_
rlabel metal2 27832 45864 27832 45864 0 _0054_
rlabel metal2 39816 33936 39816 33936 0 _0055_
rlabel metal3 35056 44520 35056 44520 0 _0056_
rlabel metal2 39592 34888 39592 34888 0 _0057_
rlabel metal2 38920 35728 38920 35728 0 _0058_
rlabel metal3 38892 31752 38892 31752 0 _0059_
rlabel metal2 41944 34776 41944 34776 0 _0060_
rlabel metal2 31360 38808 31360 38808 0 _0061_
rlabel metal3 32816 34664 32816 34664 0 _0062_
rlabel metal2 16408 39536 16408 39536 0 _0063_
rlabel metal2 3304 45752 3304 45752 0 _0064_
rlabel metal2 7336 42056 7336 42056 0 _0065_
rlabel metal2 10360 46816 10360 46816 0 _0066_
rlabel metal2 7000 45864 7000 45864 0 _0067_
rlabel metal2 10920 45813 10920 45813 0 _0068_
rlabel metal2 9688 40992 9688 40992 0 _0069_
rlabel metal2 7672 48104 7672 48104 0 _0070_
rlabel metal2 6440 44184 6440 44184 0 _0071_
rlabel metal2 13944 41720 13944 41720 0 _0072_
rlabel metal2 12824 47600 12824 47600 0 _0073_
rlabel metal2 15288 42336 15288 42336 0 _0074_
rlabel metal2 15176 40712 15176 40712 0 _0075_
rlabel metal2 7000 45304 7000 45304 0 _0076_
rlabel metal2 7000 48160 7000 48160 0 _0077_
rlabel metal2 5376 41944 5376 41944 0 _0078_
rlabel metal3 6944 45752 6944 45752 0 _0079_
rlabel via2 18088 42504 18088 42504 0 _0080_
rlabel metal2 14952 40264 14952 40264 0 _0081_
rlabel metal2 4200 45304 4200 45304 0 _0082_
rlabel metal2 6440 39256 6440 39256 0 _0083_
rlabel metal2 7112 37184 7112 37184 0 _0084_
rlabel metal2 18200 39256 18200 39256 0 _0085_
rlabel metal2 37800 34272 37800 34272 0 _0086_
rlabel metal3 20048 21672 20048 21672 0 _0087_
rlabel metal2 12936 24192 12936 24192 0 _0088_
rlabel metal3 16464 39592 16464 39592 0 _0089_
rlabel metal2 31416 39256 31416 39256 0 _0090_
rlabel metal3 34776 30184 34776 30184 0 _0091_
rlabel metal2 34328 30688 34328 30688 0 _0092_
rlabel metal2 33320 36008 33320 36008 0 _0093_
rlabel metal2 31864 38808 31864 38808 0 _0094_
rlabel metal2 4872 43568 4872 43568 0 _0095_
rlabel metal2 12264 40264 12264 40264 0 _0096_
rlabel metal2 27832 41944 27832 41944 0 _0097_
rlabel metal2 7112 40824 7112 40824 0 _0098_
rlabel metal2 7392 47320 7392 47320 0 _0099_
rlabel metal2 8680 41104 8680 41104 0 _0100_
rlabel metal2 30072 39592 30072 39592 0 _0101_
rlabel metal2 33712 39480 33712 39480 0 _0102_
rlabel metal2 32424 38780 32424 38780 0 _0103_
rlabel metal2 30744 39256 30744 39256 0 _0104_
rlabel metal3 30296 39760 30296 39760 0 _0105_
rlabel metal2 27048 42504 27048 42504 0 _0106_
rlabel metal2 16296 32256 16296 32256 0 _0107_
rlabel metal3 37464 31752 37464 31752 0 _0108_
rlabel metal2 38472 32816 38472 32816 0 _0109_
rlabel metal2 34776 39200 34776 39200 0 _0110_
rlabel metal3 33264 28056 33264 28056 0 _0111_
rlabel metal3 12040 24920 12040 24920 0 _0112_
rlabel metal3 29400 28616 29400 28616 0 _0113_
rlabel metal2 24248 28280 24248 28280 0 _0114_
rlabel metal2 39032 28840 39032 28840 0 _0115_
rlabel metal2 25368 24192 25368 24192 0 _0116_
rlabel metal3 34104 31528 34104 31528 0 _0117_
rlabel metal2 26040 28784 26040 28784 0 _0118_
rlabel via2 6888 43400 6888 43400 0 _0119_
rlabel metal3 7728 34888 7728 34888 0 _0120_
rlabel metal3 8372 23240 8372 23240 0 _0121_
rlabel metal2 29288 28672 29288 28672 0 _0122_
rlabel metal3 33152 33096 33152 33096 0 _0123_
rlabel metal2 19656 31416 19656 31416 0 _0124_
rlabel metal2 15624 24080 15624 24080 0 _0125_
rlabel metal2 28280 25984 28280 25984 0 _0126_
rlabel metal2 11704 24304 11704 24304 0 _0127_
rlabel metal3 28280 29512 28280 29512 0 _0128_
rlabel metal3 20888 39592 20888 39592 0 _0129_
rlabel metal2 21896 33544 21896 33544 0 _0130_
rlabel metal3 10752 45080 10752 45080 0 _0131_
rlabel metal2 19712 45640 19712 45640 0 _0132_
rlabel metal2 26264 34160 26264 34160 0 _0133_
rlabel via2 29064 29400 29064 29400 0 _0134_
rlabel metal2 27608 41608 27608 41608 0 _0135_
rlabel metal2 17752 32592 17752 32592 0 _0136_
rlabel metal2 19320 30408 19320 30408 0 _0137_
rlabel metal2 25032 30912 25032 30912 0 _0138_
rlabel metal2 25480 26376 25480 26376 0 _0139_
rlabel metal2 9688 34328 9688 34328 0 _0140_
rlabel metal3 19544 33208 19544 33208 0 _0141_
rlabel metal2 26320 26488 26320 26488 0 _0142_
rlabel metal2 25368 31696 25368 31696 0 _0143_
rlabel metal2 26824 32032 26824 32032 0 _0144_
rlabel metal2 17528 36904 17528 36904 0 _0145_
rlabel metal3 19152 36232 19152 36232 0 _0146_
rlabel metal2 20384 28616 20384 28616 0 _0147_
rlabel metal2 23576 29736 23576 29736 0 _0148_
rlabel metal2 24360 29288 24360 29288 0 _0149_
rlabel metal2 23968 29624 23968 29624 0 _0150_
rlabel metal2 30520 42112 30520 42112 0 _0151_
rlabel metal2 28616 42112 28616 42112 0 _0152_
rlabel metal2 13384 24080 13384 24080 0 _0153_
rlabel metal3 31024 25592 31024 25592 0 _0154_
rlabel metal2 13720 27944 13720 27944 0 _0155_
rlabel metal3 9296 43624 9296 43624 0 _0156_
rlabel metal2 8568 42392 8568 42392 0 _0157_
rlabel metal2 10248 49336 10248 49336 0 _0158_
rlabel metal2 14056 47656 14056 47656 0 _0159_
rlabel metal3 12376 43400 12376 43400 0 _0160_
rlabel metal2 16184 40600 16184 40600 0 _0161_
rlabel metal2 16520 49112 16520 49112 0 _0162_
rlabel metal3 16016 48776 16016 48776 0 _0163_
rlabel metal2 5992 42588 5992 42588 0 _0164_
rlabel metal2 5936 26264 5936 26264 0 _0165_
rlabel metal2 22904 31416 22904 31416 0 _0166_
rlabel metal2 20440 34328 20440 34328 0 _0167_
rlabel metal2 16576 40376 16576 40376 0 _0168_
rlabel metal2 16408 40880 16408 40880 0 _0169_
rlabel metal2 13720 47824 13720 47824 0 _0170_
rlabel metal2 13328 46760 13328 46760 0 _0171_
rlabel metal2 23240 25648 23240 25648 0 _0172_
rlabel metal3 19768 30184 19768 30184 0 _0173_
rlabel metal3 28504 47600 28504 47600 0 _0174_
rlabel metal2 7112 26264 7112 26264 0 _0175_
rlabel metal2 12264 41384 12264 41384 0 _0176_
rlabel metal3 28616 39872 28616 39872 0 _0177_
rlabel metal3 3220 39592 3220 39592 0 _0178_
rlabel metal3 4704 39032 4704 39032 0 _0179_
rlabel metal3 7168 30184 7168 30184 0 _0180_
rlabel metal2 6552 31304 6552 31304 0 _0181_
rlabel metal2 9016 29848 9016 29848 0 _0182_
rlabel metal2 21448 30800 21448 30800 0 _0183_
rlabel metal2 7616 25480 7616 25480 0 _0184_
rlabel metal2 7112 25816 7112 25816 0 _0185_
rlabel metal3 22456 33320 22456 33320 0 _0186_
rlabel metal2 11760 30296 11760 30296 0 _0187_
rlabel metal3 16856 35168 16856 35168 0 _0188_
rlabel metal2 19432 45528 19432 45528 0 _0189_
rlabel metal2 17640 42448 17640 42448 0 _0190_
rlabel metal2 24136 43288 24136 43288 0 _0191_
rlabel metal2 22120 44912 22120 44912 0 _0192_
rlabel metal2 18200 25984 18200 25984 0 _0193_
rlabel metal2 18032 44184 18032 44184 0 _0194_
rlabel metal3 17304 44408 17304 44408 0 _0195_
rlabel metal2 14728 24416 14728 24416 0 _0196_
rlabel metal2 23464 24864 23464 24864 0 _0197_
rlabel metal2 16072 27160 16072 27160 0 _0198_
rlabel metal2 14840 34328 14840 34328 0 _0199_
rlabel metal3 28140 25144 28140 25144 0 _0200_
rlabel metal2 15960 33600 15960 33600 0 _0201_
rlabel metal2 15848 34552 15848 34552 0 _0202_
rlabel metal2 17080 35140 17080 35140 0 _0203_
rlabel metal2 3304 34300 3304 34300 0 _0204_
rlabel metal2 2856 32984 2856 32984 0 _0205_
rlabel metal2 5432 39452 5432 39452 0 _0206_
rlabel metal2 2632 31808 2632 31808 0 _0207_
rlabel metal2 34160 39592 34160 39592 0 _0208_
rlabel metal2 30520 40768 30520 40768 0 _0209_
rlabel metal2 28840 43008 28840 43008 0 _0210_
rlabel metal2 31192 39536 31192 39536 0 _0211_
rlabel metal3 28784 38696 28784 38696 0 _0212_
rlabel metal2 7448 32256 7448 32256 0 _0213_
rlabel metal2 11816 36456 11816 36456 0 _0214_
rlabel metal2 17640 26908 17640 26908 0 _0215_
rlabel metal2 4312 31640 4312 31640 0 _0216_
rlabel metal2 2632 39200 2632 39200 0 _0217_
rlabel metal2 2464 38024 2464 38024 0 _0218_
rlabel metal2 4648 33432 4648 33432 0 _0219_
rlabel metal3 5544 33320 5544 33320 0 _0220_
rlabel metal2 14392 27160 14392 27160 0 _0221_
rlabel metal3 11536 43512 11536 43512 0 _0222_
rlabel metal3 13048 26488 13048 26488 0 _0223_
rlabel metal2 25704 27776 25704 27776 0 _0224_
rlabel metal2 24920 41216 24920 41216 0 _0225_
rlabel metal2 14056 24528 14056 24528 0 _0226_
rlabel metal2 8512 25592 8512 25592 0 _0227_
rlabel metal3 7168 28056 7168 28056 0 _0228_
rlabel metal2 16632 31584 16632 31584 0 _0229_
rlabel metal3 15428 41048 15428 41048 0 _0230_
rlabel metal2 18200 41608 18200 41608 0 _0231_
rlabel metal2 18648 24752 18648 24752 0 _0232_
rlabel metal2 19208 22904 19208 22904 0 _0233_
rlabel metal3 17304 24696 17304 24696 0 _0234_
rlabel metal3 23800 24808 23800 24808 0 _0235_
rlabel metal2 18648 44408 18648 44408 0 _0236_
rlabel metal2 9912 24640 9912 24640 0 _0237_
rlabel metal2 21112 24248 21112 24248 0 _0238_
rlabel metal2 14224 26488 14224 26488 0 _0239_
rlabel metal2 20440 25088 20440 25088 0 _0240_
rlabel metal2 19096 26376 19096 26376 0 _0241_
rlabel metal2 18312 32984 18312 32984 0 _0242_
rlabel metal2 22792 25760 22792 25760 0 _0243_
rlabel metal2 20888 36176 20888 36176 0 _0244_
rlabel metal2 20776 33656 20776 33656 0 _0245_
rlabel metal2 23016 35168 23016 35168 0 _0246_
rlabel metal2 8792 25480 8792 25480 0 _0247_
rlabel metal2 22008 25256 22008 25256 0 _0248_
rlabel metal2 7728 37240 7728 37240 0 _0249_
rlabel metal2 19992 38668 19992 38668 0 _0250_
rlabel metal2 25816 36736 25816 36736 0 _0251_
rlabel metal2 23912 36008 23912 36008 0 _0252_
rlabel metal2 23240 36792 23240 36792 0 _0253_
rlabel metal2 15512 30408 15512 30408 0 _0254_
rlabel metal2 20048 35448 20048 35448 0 _0255_
rlabel metal2 21000 34496 21000 34496 0 _0256_
rlabel metal2 20160 35672 20160 35672 0 _0257_
rlabel metal2 18984 37912 18984 37912 0 _0258_
rlabel metal2 17192 31640 17192 31640 0 _0259_
rlabel metal2 19096 34048 19096 34048 0 _0260_
rlabel metal3 22008 34328 22008 34328 0 _0261_
rlabel metal2 24696 36568 24696 36568 0 _0262_
rlabel metal2 25256 37968 25256 37968 0 _0263_
rlabel metal2 26936 43176 26936 43176 0 _0264_
rlabel metal3 10024 39032 10024 39032 0 _0265_
rlabel metal2 16072 29120 16072 29120 0 _0266_
rlabel metal3 22624 27048 22624 27048 0 _0267_
rlabel metal2 24640 30968 24640 30968 0 _0268_
rlabel metal2 26040 31808 26040 31808 0 _0269_
rlabel metal3 19656 37576 19656 37576 0 _0270_
rlabel metal2 10248 25760 10248 25760 0 _0271_
rlabel metal3 9296 25480 9296 25480 0 _0272_
rlabel metal2 10472 25424 10472 25424 0 _0273_
rlabel metal3 11704 25368 11704 25368 0 _0274_
rlabel metal3 11648 25256 11648 25256 0 _0275_
rlabel metal2 11928 47208 11928 47208 0 _0276_
rlabel metal2 11816 26152 11816 26152 0 _0277_
rlabel metal3 11480 25480 11480 25480 0 _0278_
rlabel metal2 11368 24416 11368 24416 0 _0279_
rlabel metal2 28280 43120 28280 43120 0 _0280_
rlabel metal2 26040 45920 26040 45920 0 _0281_
rlabel metal3 27832 48216 27832 48216 0 _0282_
rlabel metal2 28728 43568 28728 43568 0 _0283_
rlabel metal2 29848 44380 29848 44380 0 _0284_
rlabel metal2 16128 46648 16128 46648 0 _0285_
rlabel metal2 15960 47040 15960 47040 0 _0286_
rlabel metal2 23184 41832 23184 41832 0 _0287_
rlabel metal2 17024 45864 17024 45864 0 _0288_
rlabel metal2 16128 44408 16128 44408 0 _0289_
rlabel metal2 19768 45136 19768 45136 0 _0290_
rlabel metal3 17304 47432 17304 47432 0 _0291_
rlabel metal2 17416 45416 17416 45416 0 _0292_
rlabel metal2 18536 32536 18536 32536 0 _0293_
rlabel metal2 15512 41160 15512 41160 0 _0294_
rlabel metal2 17528 41776 17528 41776 0 _0295_
rlabel metal2 16408 44016 16408 44016 0 _0296_
rlabel metal2 2296 31528 2296 31528 0 _0297_
rlabel metal3 6328 35896 6328 35896 0 _0298_
rlabel metal2 4088 34496 4088 34496 0 _0299_
rlabel metal2 16632 44128 16632 44128 0 _0300_
rlabel metal2 18088 31304 18088 31304 0 _0301_
rlabel metal3 13048 34888 13048 34888 0 _0302_
rlabel metal2 17864 31360 17864 31360 0 _0303_
rlabel metal2 16296 30800 16296 30800 0 _0304_
rlabel metal2 17976 42000 17976 42000 0 _0305_
rlabel metal2 16688 39816 16688 39816 0 _0306_
rlabel metal3 17472 44296 17472 44296 0 _0307_
rlabel metal2 17304 44800 17304 44800 0 _0308_
rlabel metal2 30072 37184 30072 37184 0 _0309_
rlabel metal2 29792 37464 29792 37464 0 _0310_
rlabel metal2 28728 37184 28728 37184 0 _0311_
rlabel metal3 26880 38920 26880 38920 0 _0312_
rlabel metal2 28616 41384 28616 41384 0 _0313_
rlabel metal2 25816 40376 25816 40376 0 _0314_
rlabel metal2 25144 32480 25144 32480 0 _0315_
rlabel metal2 23016 25368 23016 25368 0 _0316_
rlabel metal2 25816 38080 25816 38080 0 _0317_
rlabel metal2 12376 36456 12376 36456 0 _0318_
rlabel metal2 28056 37968 28056 37968 0 _0319_
rlabel metal3 19992 38136 19992 38136 0 _0320_
rlabel metal2 20552 40992 20552 40992 0 _0321_
rlabel metal3 22960 38696 22960 38696 0 _0322_
rlabel metal2 25144 41216 25144 41216 0 _0323_
rlabel metal2 27384 47488 27384 47488 0 _0324_
rlabel metal3 25928 49000 25928 49000 0 _0325_
rlabel metal3 24248 33432 24248 33432 0 _0326_
rlabel metal2 28392 38864 28392 38864 0 _0327_
rlabel metal3 28504 34664 28504 34664 0 _0328_
rlabel metal3 28728 34216 28728 34216 0 _0329_
rlabel metal2 28392 39592 28392 39592 0 _0330_
rlabel metal2 28000 38920 28000 38920 0 _0331_
rlabel metal2 2912 34776 2912 34776 0 _0332_
rlabel metal2 18200 40712 18200 40712 0 _0333_
rlabel metal3 15316 27832 15316 27832 0 _0334_
rlabel metal2 18704 37240 18704 37240 0 _0335_
rlabel metal2 19096 36400 19096 36400 0 _0336_
rlabel metal2 19320 34944 19320 34944 0 _0337_
rlabel metal2 17416 37464 17416 37464 0 _0338_
rlabel metal2 17640 34048 17640 34048 0 _0339_
rlabel metal2 16296 37296 16296 37296 0 _0340_
rlabel metal3 18256 38024 18256 38024 0 _0341_
rlabel metal3 20944 30072 20944 30072 0 _0342_
rlabel metal3 19096 28616 19096 28616 0 _0343_
rlabel metal2 18200 28336 18200 28336 0 _0344_
rlabel metal3 18592 23240 18592 23240 0 _0345_
rlabel metal2 18872 26992 18872 26992 0 _0346_
rlabel metal2 18424 27160 18424 27160 0 _0347_
rlabel metal3 10584 26488 10584 26488 0 _0348_
rlabel metal2 9800 26656 9800 26656 0 _0349_
rlabel metal2 17752 27160 17752 27160 0 _0350_
rlabel metal3 18144 30968 18144 30968 0 _0351_
rlabel metal2 18816 39032 18816 39032 0 _0352_
rlabel metal2 17864 42392 17864 42392 0 _0353_
rlabel metal2 20328 41888 20328 41888 0 _0354_
rlabel metal2 19656 41272 19656 41272 0 _0355_
rlabel metal2 18648 48776 18648 48776 0 _0356_
rlabel metal2 18704 41944 18704 41944 0 _0357_
rlabel metal2 18368 41832 18368 41832 0 _0358_
rlabel metal3 19152 40376 19152 40376 0 _0359_
rlabel metal2 19544 41104 19544 41104 0 _0360_
rlabel metal3 25984 45752 25984 45752 0 _0361_
rlabel metal3 28728 37128 28728 37128 0 _0362_
rlabel metal2 27384 35112 27384 35112 0 _0363_
rlabel metal2 27832 32088 27832 32088 0 _0364_
rlabel metal3 22596 31864 22596 31864 0 _0365_
rlabel metal2 27776 31192 27776 31192 0 _0366_
rlabel metal2 27328 43512 27328 43512 0 _0367_
rlabel metal2 26824 45136 26824 45136 0 _0368_
rlabel metal2 5544 26572 5544 26572 0 _0369_
rlabel metal2 8904 33376 8904 33376 0 _0370_
rlabel metal2 10752 29960 10752 29960 0 _0371_
rlabel metal2 29176 41216 29176 41216 0 _0372_
rlabel metal3 14168 29400 14168 29400 0 _0373_
rlabel metal2 15064 28784 15064 28784 0 _0374_
rlabel metal2 14728 29848 14728 29848 0 _0375_
rlabel metal2 23800 40712 23800 40712 0 _0376_
rlabel metal2 24808 45136 24808 45136 0 _0377_
rlabel metal2 22400 48104 22400 48104 0 _0378_
rlabel metal2 21896 48160 21896 48160 0 _0379_
rlabel metal2 23912 48384 23912 48384 0 _0380_
rlabel metal2 24024 47152 24024 47152 0 _0381_
rlabel metal2 26936 46760 26936 46760 0 _0382_
rlabel metal2 27720 48496 27720 48496 0 _0383_
rlabel metal2 28392 43232 28392 43232 0 _0384_
rlabel metal2 27160 43288 27160 43288 0 _0385_
rlabel metal2 29624 45584 29624 45584 0 _0386_
rlabel metal2 25368 41888 25368 41888 0 _0387_
rlabel metal2 25816 28616 25816 28616 0 _0388_
rlabel metal2 26376 30520 26376 30520 0 _0389_
rlabel metal2 26600 30520 26600 30520 0 _0390_
rlabel metal2 26040 40152 26040 40152 0 _0391_
rlabel metal2 25648 40600 25648 40600 0 _0392_
rlabel metal3 20440 28616 20440 28616 0 _0393_
rlabel metal2 10080 36680 10080 36680 0 _0394_
rlabel metal2 8680 28784 8680 28784 0 _0395_
rlabel metal2 10696 29064 10696 29064 0 _0396_
rlabel metal2 10136 28896 10136 28896 0 _0397_
rlabel metal2 5712 31080 5712 31080 0 _0398_
rlabel metal2 3416 30968 3416 30968 0 _0399_
rlabel metal2 6328 29736 6328 29736 0 _0400_
rlabel metal2 2520 41552 2520 41552 0 _0401_
rlabel metal3 2352 44856 2352 44856 0 _0402_
rlabel metal2 14056 25424 14056 25424 0 _0403_
rlabel metal2 10304 26376 10304 26376 0 _0404_
rlabel metal3 7952 27160 7952 27160 0 _0405_
rlabel metal3 7840 26488 7840 26488 0 _0406_
rlabel metal2 5320 27776 5320 27776 0 _0407_
rlabel metal2 7112 28280 7112 28280 0 _0408_
rlabel metal2 23128 43288 23128 43288 0 _0409_
rlabel metal2 20664 40544 20664 40544 0 _0410_
rlabel metal2 21504 39032 21504 39032 0 _0411_
rlabel metal3 23016 48104 23016 48104 0 _0412_
rlabel metal3 18760 48888 18760 48888 0 _0413_
rlabel metal2 19992 49056 19992 49056 0 _0414_
rlabel metal2 25928 44352 25928 44352 0 _0415_
rlabel metal2 29176 46256 29176 46256 0 _0416_
rlabel metal2 38696 46144 38696 46144 0 _0417_
rlabel metal3 30464 44520 30464 44520 0 _0418_
rlabel metal2 20328 47712 20328 47712 0 _0419_
rlabel metal2 22008 44856 22008 44856 0 _0420_
rlabel metal2 22792 45360 22792 45360 0 _0421_
rlabel metal2 19656 28952 19656 28952 0 _0422_
rlabel metal2 18760 35336 18760 35336 0 _0423_
rlabel metal3 16128 26376 16128 26376 0 _0424_
rlabel metal2 17528 35672 17528 35672 0 _0425_
rlabel metal2 3752 27216 3752 27216 0 _0426_
rlabel metal2 3192 42728 3192 42728 0 _0427_
rlabel metal2 2912 35000 2912 35000 0 _0428_
rlabel metal2 17752 35616 17752 35616 0 _0429_
rlabel metal2 22736 40040 22736 40040 0 _0430_
rlabel metal2 29400 45584 29400 45584 0 _0431_
rlabel metal2 26376 33544 26376 33544 0 _0432_
rlabel metal2 30240 41944 30240 41944 0 _0433_
rlabel metal3 29176 42728 29176 42728 0 _0434_
rlabel metal2 29288 43960 29288 43960 0 _0435_
rlabel metal2 33880 41440 33880 41440 0 _0436_
rlabel metal3 27440 38696 27440 38696 0 _0437_
rlabel metal2 26936 40320 26936 40320 0 _0438_
rlabel metal3 20160 39032 20160 39032 0 _0439_
rlabel metal2 20440 37240 20440 37240 0 _0440_
rlabel metal2 21560 38724 21560 38724 0 _0441_
rlabel metal3 26040 38920 26040 38920 0 _0442_
rlabel metal3 13104 38808 13104 38808 0 _0443_
rlabel metal2 9240 31416 9240 31416 0 _0444_
rlabel metal2 3640 36904 3640 36904 0 _0445_
rlabel metal2 28168 48720 28168 48720 0 _0446_
rlabel metal2 27608 40096 27608 40096 0 _0447_
rlabel metal2 20720 24136 20720 24136 0 _0448_
rlabel metal2 15288 27272 15288 27272 0 _0449_
rlabel metal2 15848 27720 15848 27720 0 _0450_
rlabel metal2 31696 39816 31696 39816 0 _0451_
rlabel metal2 27048 39480 27048 39480 0 _0452_
rlabel metal2 17640 25256 17640 25256 0 _0453_
rlabel metal2 16184 23408 16184 23408 0 _0454_
rlabel metal2 16576 25592 16576 25592 0 _0455_
rlabel metal3 20664 24024 20664 24024 0 _0456_
rlabel metal2 23240 48216 23240 48216 0 _0457_
rlabel metal2 23744 48216 23744 48216 0 _0458_
rlabel metal2 26824 40712 26824 40712 0 _0459_
rlabel metal2 33544 43008 33544 43008 0 _0460_
rlabel metal2 30408 43064 30408 43064 0 _0461_
rlabel metal2 31080 43008 31080 43008 0 _0462_
rlabel metal2 21560 41384 21560 41384 0 _0463_
rlabel metal2 19600 39928 19600 39928 0 _0464_
rlabel metal2 21560 30688 21560 30688 0 _0465_
rlabel metal3 20720 29624 20720 29624 0 _0466_
rlabel metal2 21840 30408 21840 30408 0 _0467_
rlabel metal2 22120 41664 22120 41664 0 _0468_
rlabel metal3 9464 38584 9464 38584 0 _0469_
rlabel metal2 2968 40544 2968 40544 0 _0470_
rlabel metal2 4256 36456 4256 36456 0 _0471_
rlabel metal2 8232 37744 8232 37744 0 _0472_
rlabel metal2 21560 41776 21560 41776 0 _0473_
rlabel metal3 20720 46648 20720 46648 0 _0474_
rlabel metal2 21392 45304 21392 45304 0 _0475_
rlabel metal2 22456 43680 22456 43680 0 _0476_
rlabel metal2 30968 42224 30968 42224 0 _0477_
rlabel metal3 35336 43512 35336 43512 0 _0478_
rlabel metal2 28728 39984 28728 39984 0 _0479_
rlabel metal2 30800 42728 30800 42728 0 _0480_
rlabel metal2 19208 48720 19208 48720 0 _0481_
rlabel metal2 20104 48328 20104 48328 0 _0482_
rlabel metal2 19992 47824 19992 47824 0 _0483_
rlabel metal2 12936 30296 12936 30296 0 _0484_
rlabel metal3 14560 36680 14560 36680 0 _0485_
rlabel metal2 15064 36568 15064 36568 0 _0486_
rlabel metal3 15680 37016 15680 37016 0 _0487_
rlabel metal2 15344 38584 15344 38584 0 _0488_
rlabel metal3 17248 43512 17248 43512 0 _0489_
rlabel metal2 2856 43008 2856 43008 0 _0490_
rlabel metal2 2632 30184 2632 30184 0 _0491_
rlabel metal2 18648 43008 18648 43008 0 _0492_
rlabel metal2 30632 44072 30632 44072 0 _0493_
rlabel metal3 29456 54488 29456 54488 0 _0494_
rlabel metal3 10248 52920 10248 52920 0 _0495_
rlabel metal2 12488 54432 12488 54432 0 _0496_
rlabel metal2 13832 53984 13832 53984 0 _0497_
rlabel via2 11704 52696 11704 52696 0 _0498_
rlabel metal2 30296 47376 30296 47376 0 _0499_
rlabel metal2 11256 50876 11256 50876 0 _0500_
rlabel metal2 29176 53312 29176 53312 0 _0501_
rlabel metal3 11200 51576 11200 51576 0 _0502_
rlabel metal3 11256 53480 11256 53480 0 _0503_
rlabel metal2 11424 50456 11424 50456 0 _0504_
rlabel metal2 29512 52360 29512 52360 0 _0505_
rlabel metal3 33040 41944 33040 41944 0 _0506_
rlabel metal2 12096 52136 12096 52136 0 _0507_
rlabel metal2 32648 49672 32648 49672 0 _0508_
rlabel metal3 34216 43624 34216 43624 0 _0509_
rlabel metal2 34552 44912 34552 44912 0 _0510_
rlabel metal2 36120 41608 36120 41608 0 _0511_
rlabel metal2 36064 48776 36064 48776 0 _0512_
rlabel metal2 34664 40712 34664 40712 0 _0513_
rlabel metal2 41272 52360 41272 52360 0 _0514_
rlabel metal3 35168 40376 35168 40376 0 _0515_
rlabel metal3 40768 54376 40768 54376 0 _0516_
rlabel metal2 34216 45136 34216 45136 0 _0517_
rlabel metal2 38472 49504 38472 49504 0 _0518_
rlabel metal3 24528 50232 24528 50232 0 _0519_
rlabel metal2 26264 52752 26264 52752 0 _0520_
rlabel metal2 27552 52808 27552 52808 0 _0521_
rlabel metal2 25424 52920 25424 52920 0 _0522_
rlabel metal3 23968 50456 23968 50456 0 _0523_
rlabel metal3 25760 53816 25760 53816 0 _0524_
rlabel metal3 23296 53816 23296 53816 0 _0525_
rlabel metal3 26432 50568 26432 50568 0 _0526_
rlabel metal2 39032 45528 39032 45528 0 _0527_
rlabel metal2 39480 46648 39480 46648 0 _0528_
rlabel metal2 38864 47208 38864 47208 0 _0529_
rlabel metal3 40264 46760 40264 46760 0 _0530_
rlabel metal2 41048 43064 41048 43064 0 _0531_
rlabel metal2 39592 44408 39592 44408 0 _0532_
rlabel metal2 41160 45080 41160 45080 0 _0533_
rlabel metal2 29848 53760 29848 53760 0 _0534_
rlabel metal2 30408 54040 30408 54040 0 _0535_
rlabel metal2 31864 53872 31864 53872 0 _0536_
rlabel metal2 31752 54432 31752 54432 0 _0537_
rlabel metal2 31864 52864 31864 52864 0 _0538_
rlabel metal2 33992 54432 33992 54432 0 _0539_
rlabel metal2 42280 52528 42280 52528 0 _0540_
rlabel metal2 37128 52584 37128 52584 0 _0541_
rlabel metal3 40264 54600 40264 54600 0 _0542_
rlabel metal3 40152 54488 40152 54488 0 _0543_
rlabel metal2 39256 51352 39256 51352 0 _0544_
rlabel metal2 41720 53368 41720 53368 0 _0545_
rlabel metal2 41832 51296 41832 51296 0 _0546_
rlabel metal2 41384 53928 41384 53928 0 _0547_
rlabel metal2 30296 50680 30296 50680 0 _0548_
rlabel metal2 14616 53312 14616 53312 0 _0549_
rlabel metal3 16184 51912 16184 51912 0 _0550_
rlabel metal2 18872 52528 18872 52528 0 _0551_
rlabel metal2 15176 54656 15176 54656 0 _0552_
rlabel metal2 15176 52248 15176 52248 0 _0553_
rlabel metal3 18144 54488 18144 54488 0 _0554_
rlabel metal2 18312 51408 18312 51408 0 _0555_
rlabel metal2 31192 47936 31192 47936 0 _0556_
rlabel metal2 30632 49728 30632 49728 0 _0557_
rlabel metal3 33992 48776 33992 48776 0 _0558_
rlabel metal2 32872 46312 32872 46312 0 _0559_
rlabel metal3 34720 49000 34720 49000 0 _0560_
rlabel metal2 34440 46648 34440 46648 0 _0561_
rlabel metal2 31864 48552 31864 48552 0 _0562_
rlabel metal2 23128 57778 23128 57778 0 bus_in[0]
rlabel metal2 25368 57778 25368 57778 0 bus_in[1]
rlabel metal2 27944 55888 27944 55888 0 bus_in[2]
rlabel metal2 29848 57778 29848 57778 0 bus_in[3]
rlabel metal2 32088 57778 32088 57778 0 bus_in[4]
rlabel metal2 34328 57778 34328 57778 0 bus_in[5]
rlabel metal2 36568 57778 36568 57778 0 bus_in[6]
rlabel metal2 39368 56448 39368 56448 0 bus_in[7]
rlabel metal2 41048 57778 41048 57778 0 bus_out[0]
rlabel metal2 43288 57778 43288 57778 0 bus_out[1]
rlabel metal3 46144 55384 46144 55384 0 bus_out[2]
rlabel metal2 47768 57778 47768 57778 0 bus_out[3]
rlabel metal2 50008 57778 50008 57778 0 bus_out[4]
rlabel metal3 53032 55384 53032 55384 0 bus_out[5]
rlabel metal2 54488 57778 54488 57778 0 bus_out[6]
rlabel metal2 56728 57330 56728 57330 0 bus_out[7]
rlabel metal2 30184 46872 30184 46872 0 clknet_0_wb_clk_i
rlabel metal2 20776 53312 20776 53312 0 clknet_2_0__leaf_wb_clk_i
rlabel metal3 6048 51352 6048 51352 0 clknet_2_1__leaf_wb_clk_i
rlabel metal3 35560 43736 35560 43736 0 clknet_2_2__leaf_wb_clk_i
rlabel metal3 41272 48104 41272 48104 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 16464 56280 16464 56280 0 cs_port[0]
rlabel metal2 18648 57778 18648 57778 0 cs_port[1]
rlabel metal2 21000 56168 21000 56168 0 cs_port[2]
rlabel metal2 2184 48552 2184 48552 0 full_addr\[0\]
rlabel metal2 36456 53648 36456 53648 0 full_addr\[10\]
rlabel metal3 36624 52248 36624 52248 0 full_addr\[11\]
rlabel metal2 40320 51464 40320 51464 0 full_addr\[12\]
rlabel metal2 42616 52920 42616 52920 0 full_addr\[13\]
rlabel metal2 42504 50904 42504 50904 0 full_addr\[14\]
rlabel metal2 42952 53760 42952 53760 0 full_addr\[15\]
rlabel metal2 2184 50680 2184 50680 0 full_addr\[1\]
rlabel metal3 6608 50792 6608 50792 0 full_addr\[2\]
rlabel metal2 7112 50960 7112 50960 0 full_addr\[3\]
rlabel metal3 38864 38696 38864 38696 0 full_addr\[4\]
rlabel metal2 38696 35000 38696 35000 0 full_addr\[5\]
rlabel metal2 40376 38024 40376 38024 0 full_addr\[6\]
rlabel metal3 37632 40488 37632 40488 0 full_addr\[7\]
rlabel metal2 32088 53984 32088 53984 0 full_addr\[8\]
rlabel metal3 34384 53032 34384 53032 0 full_addr\[9\]
rlabel metal2 11928 57778 11928 57778 0 le_hi_act
rlabel metal2 9688 57778 9688 57778 0 le_lo_act
rlabel metal2 8120 55440 8120 55440 0 net1
rlabel metal2 18088 49056 18088 49056 0 net10
rlabel metal2 18312 48552 18312 48552 0 net11
rlabel metal3 20776 45864 20776 45864 0 net12
rlabel metal2 29288 54208 29288 54208 0 net13
rlabel metal2 28616 48720 28616 48720 0 net14
rlabel metal2 2072 30184 2072 30184 0 net15
rlabel metal2 1960 48776 1960 48776 0 net16
rlabel metal2 2800 51464 2800 51464 0 net17
rlabel metal1 2464 52696 2464 52696 0 net18
rlabel metal3 1848 54600 1848 54600 0 net19
rlabel metal2 23016 55496 23016 55496 0 net2
rlabel metal2 2016 55440 2016 55440 0 net20
rlabel metal2 2408 49840 2408 49840 0 net21
rlabel metal3 2968 33096 2968 33096 0 net22
rlabel metal2 6440 33376 6440 33376 0 net23
rlabel metal3 2464 31080 2464 31080 0 net24
rlabel metal2 2744 35056 2744 35056 0 net25
rlabel metal3 1568 39592 1568 39592 0 net26
rlabel metal2 2072 41496 2072 41496 0 net27
rlabel metal2 2072 43064 2072 43064 0 net28
rlabel metal2 2632 38276 2632 38276 0 net29
rlabel metal2 25536 55272 25536 55272 0 net3
rlabel metal2 2240 35784 2240 35784 0 net30
rlabel metal2 2352 3640 2352 3640 0 net31
rlabel metal2 2072 21224 2072 21224 0 net32
rlabel metal2 2128 22232 2128 22232 0 net33
rlabel metal4 2072 29288 2072 29288 0 net34
rlabel metal3 2352 36008 2352 36008 0 net35
rlabel metal2 2072 28280 2072 28280 0 net36
rlabel metal2 2800 28616 2800 28616 0 net37
rlabel metal2 1848 4536 1848 4536 0 net38
rlabel metal2 2184 5824 2184 5824 0 net39
rlabel metal2 28056 56168 28056 56168 0 net4
rlabel metal3 3864 9464 3864 9464 0 net40
rlabel metal3 5264 26824 5264 26824 0 net41
rlabel metal2 2016 11256 2016 11256 0 net42
rlabel metal2 2072 13104 2072 13104 0 net43
rlabel metal2 2520 21112 2520 21112 0 net44
rlabel metal2 2128 20440 2128 20440 0 net45
rlabel metal3 1512 23464 1512 23464 0 net46
rlabel metal2 13720 54964 13720 54964 0 net47
rlabel metal2 5880 55664 5880 55664 0 net48
rlabel metal2 28280 49280 28280 49280 0 net49
rlabel metal2 29624 53592 29624 53592 0 net5
rlabel metal2 43736 55552 43736 55552 0 net50
rlabel metal2 45416 52024 45416 52024 0 net51
rlabel metal2 47880 56056 47880 56056 0 net52
rlabel metal2 50904 54432 50904 54432 0 net53
rlabel metal2 52416 55048 52416 55048 0 net54
rlabel metal3 49616 53816 49616 53816 0 net55
rlabel metal2 55384 49392 55384 49392 0 net56
rlabel metal2 32648 55720 32648 55720 0 net6
rlabel metal2 34888 55328 34888 55328 0 net7
rlabel metal2 37128 55720 37128 55720 0 net8
rlabel metal2 39144 55412 39144 55412 0 net9
rlabel metal2 1736 30464 1736 30464 0 ram_end[0]
rlabel metal2 1736 48776 1736 48776 0 ram_end[10]
rlabel metal2 1848 50904 1848 50904 0 ram_end[11]
rlabel metal2 1736 52584 1736 52584 0 ram_end[12]
rlabel metal2 1736 54264 1736 54264 0 ram_end[13]
rlabel metal2 1736 55944 1736 55944 0 ram_end[14]
rlabel metal3 1470 57624 1470 57624 0 ram_end[15]
rlabel metal2 1736 32872 1736 32872 0 ram_end[1]
rlabel metal3 1246 34328 1246 34328 0 ram_end[2]
rlabel metal2 1736 36680 1736 36680 0 ram_end[3]
rlabel metal2 1848 38668 1848 38668 0 ram_end[4]
rlabel metal2 1736 40040 1736 40040 0 ram_end[5]
rlabel metal2 1736 41328 1736 41328 0 ram_end[6]
rlabel metal2 1848 43344 1848 43344 0 ram_end[7]
rlabel metal2 1736 45416 1736 45416 0 ram_end[8]
rlabel metal2 1736 46816 1736 46816 0 ram_end[9]
rlabel metal2 1736 2744 1736 2744 0 ram_start[0]
rlabel metal3 1246 19992 1246 19992 0 ram_start[10]
rlabel metal2 1736 22008 1736 22008 0 ram_start[11]
rlabel metal2 1736 23688 1736 23688 0 ram_start[12]
rlabel metal3 1246 25368 1246 25368 0 ram_start[13]
rlabel metal2 1736 27496 1736 27496 0 ram_start[14]
rlabel metal2 2408 29512 2408 29512 0 ram_start[15]
rlabel metal2 1736 4088 1736 4088 0 ram_start[1]
rlabel metal2 1736 5768 1736 5768 0 ram_start[2]
rlabel metal2 1736 7784 1736 7784 0 ram_start[3]
rlabel metal2 1736 9464 1736 9464 0 ram_start[4]
rlabel metal2 1736 11144 1736 11144 0 ram_start[5]
rlabel metal3 1246 12824 1246 12824 0 ram_start[6]
rlabel metal2 1736 14952 1736 14952 0 ram_start[7]
rlabel metal2 1736 16632 1736 16632 0 ram_start[8]
rlabel metal2 1736 18312 1736 18312 0 ram_start[9]
rlabel metal2 14168 57778 14168 57778 0 rom_enabled
rlabel metal2 5152 56280 5152 56280 0 rst
rlabel metal3 4312 53816 4312 53816 0 wb_clk_i
rlabel metal2 24528 50120 24528 50120 0 writable\[0\]
rlabel metal2 23016 49224 23016 49224 0 writable\[10\]
rlabel metal3 20328 49896 20328 49896 0 writable\[11\]
rlabel metal2 29568 49112 29568 49112 0 writable\[12\]
rlabel metal2 34384 48776 34384 48776 0 writable\[13\]
rlabel metal2 34552 46200 34552 46200 0 writable\[14\]
rlabel metal2 29288 49280 29288 49280 0 writable\[15\]
rlabel metal2 28168 54096 28168 54096 0 writable\[1\]
rlabel metal2 24584 49392 24584 49392 0 writable\[2\]
rlabel metal2 27608 50568 27608 50568 0 writable\[3\]
rlabel metal2 39480 47096 39480 47096 0 writable\[4\]
rlabel metal2 41384 42728 41384 42728 0 writable\[5\]
rlabel metal3 38024 43624 38024 43624 0 writable\[6\]
rlabel metal2 41048 44632 41048 44632 0 writable\[7\]
rlabel metal2 16408 49644 16408 49644 0 writable\[8\]
rlabel metal2 16072 51296 16072 51296 0 writable\[9\]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
