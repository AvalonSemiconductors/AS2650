* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

.subckt wrapped_as2650 RAM_end_addr[0] RAM_end_addr[10] RAM_end_addr[11] RAM_end_addr[12]
+ RAM_end_addr[13] RAM_end_addr[14] RAM_end_addr[15] RAM_end_addr[1] RAM_end_addr[2]
+ RAM_end_addr[3] RAM_end_addr[4] RAM_end_addr[5] RAM_end_addr[6] RAM_end_addr[7]
+ RAM_end_addr[8] RAM_end_addr[9] RAM_start_addr[0] RAM_start_addr[10] RAM_start_addr[11]
+ RAM_start_addr[12] RAM_start_addr[13] RAM_start_addr[14] RAM_start_addr[15] RAM_start_addr[1]
+ RAM_start_addr[2] RAM_start_addr[3] RAM_start_addr[4] RAM_start_addr[5] RAM_start_addr[6]
+ RAM_start_addr[7] RAM_start_addr[8] RAM_start_addr[9] WEb_ram boot_rom_en bus_addr[0]
+ bus_addr[1] bus_addr[2] bus_addr[3] bus_addr[4] bus_addr[5] bus_cyc bus_data_out[0]
+ bus_data_out[1] bus_data_out[2] bus_data_out[3] bus_data_out[4] bus_data_out[5]
+ bus_data_out[6] bus_data_out[7] bus_in_gpios[0] bus_in_gpios[1] bus_in_gpios[2]
+ bus_in_gpios[3] bus_in_gpios[4] bus_in_gpios[5] bus_in_gpios[6] bus_in_gpios[7]
+ bus_in_serial_ports[0] bus_in_serial_ports[1] bus_in_serial_ports[2] bus_in_serial_ports[3]
+ bus_in_serial_ports[4] bus_in_serial_ports[5] bus_in_serial_ports[6] bus_in_serial_ports[7]
+ bus_in_sid[0] bus_in_sid[1] bus_in_sid[2] bus_in_sid[3] bus_in_sid[4] bus_in_sid[5]
+ bus_in_sid[6] bus_in_sid[7] bus_in_timers[0] bus_in_timers[1] bus_in_timers[2] bus_in_timers[3]
+ bus_in_timers[4] bus_in_timers[5] bus_in_timers[6] bus_in_timers[7] bus_we_gpios
+ bus_we_serial_ports bus_we_sid bus_we_timers cs_port[0] cs_port[1] cs_port[2] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8]
+ io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[1] io_out[2]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1]
+ irq[2] irqs[0] irqs[1] irqs[2] irqs[3] irqs[4] irqs[5] irqs[6] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] last_addr[0] last_addr[10] last_addr[11] last_addr[12] last_addr[13]
+ last_addr[14] last_addr[15] last_addr[1] last_addr[2] last_addr[3] last_addr[4]
+ last_addr[5] last_addr[6] last_addr[7] last_addr[8] last_addr[9] le_hi_act le_lo_act
+ ram_bus_in[0] ram_bus_in[1] ram_bus_in[2] ram_bus_in[3] ram_bus_in[4] ram_bus_in[5]
+ ram_bus_in[6] ram_bus_in[7] ram_enabled requested_addr[0] requested_addr[10] requested_addr[11]
+ requested_addr[12] requested_addr[13] requested_addr[14] requested_addr[15] requested_addr[1]
+ requested_addr[2] requested_addr[3] requested_addr[4] requested_addr[5] requested_addr[6]
+ requested_addr[7] requested_addr[8] requested_addr[9] reset_out rom_bus_in[0] rom_bus_in[1]
+ rom_bus_in[2] rom_bus_in[3] rom_bus_in[4] rom_bus_in[5] rom_bus_in[6] rom_bus_in[7]
+ rom_bus_out[0] rom_bus_out[1] rom_bus_out[2] rom_bus_out[3] rom_bus_out[4] rom_bus_out[5]
+ rom_bus_out[6] rom_bus_out[7] vdd vss wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i wbs_we_i la_data_out[39] la_data_out[38]
+ la_data_out[55]
XFILLER_0_78_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05903_ _00796_ as2650.regs\[7\]\[4\] _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09671_ _03745_ _02814_ _02790_ _03857_ _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06883_ _01800_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05834_ _00707_ as2650.regs\[7\]\[0\] _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08622_ _03058_ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_307 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_318 irq[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_329 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_08553_ as2650.stack\[4\]\[1\] _03249_ _03251_ as2650.stack\[5\]\[1\] _03256_ _03257_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_49_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05765_ _00768_ _00775_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07137__I1 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07504_ net182 _02060_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08484_ _03186_ _03188_ _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05696_ as2650.regs\[2\]\[7\] _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07435_ _02192_ _01950_ _02262_ _02148_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_4_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08942__I _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07366_ _02181_ wb_counter\[13\] _02203_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06317_ _01275_ _01287_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09105_ _01771_ _02616_ _03794_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08262__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07297_ _02116_ _02140_ _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08163__B _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07558__I _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06273__A1 _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09036_ _03727_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06248_ _01128_ _01220_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_148_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_148_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06179_ _01142_ _01151_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_143_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09938_ _01465_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05806__I _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09869_ as2650.stack\[5\]\[4\] _04534_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_1543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05742__S _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09278__A1 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07128__I1 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_104_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11085__A1 _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11762_ _00541_ clknet_leaf_5_wb_clk_i as2650.stack\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_120_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10713_ as2650.stack\[8\]\[2\] _05191_ _05194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_137_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11693_ _00477_ clknet_leaf_79_wb_clk_i as2650.regs\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10644_ _05150_ _05151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10575_ as2650.stack\[15\]\[11\] _05096_ _05103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer7 _01072_ net351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06372__I _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07461__B1 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10060__A2 _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_90_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_2_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09753__A2 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08299__I _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07417__B _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ as2650.stack\[14\]\[12\] _05515_ _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05716__I _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_143_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11058_ as2650.stack\[0\]\[12\] _05471_ _05472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_88_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_60_wb_clk_i clknet_4_12__leaf_wb_clk_i clknet_leaf_60_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10009_ _01959_ _04615_ _04620_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_47_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10823__A1 _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07220_ _02072_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09858__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07151_ net409 _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06102_ _01078_ net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06282__I _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold103_I wbs_dat_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06255__A1 _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07082_ _01820_ _01980_ _01982_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06033_ _01021_ net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_2_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11000__A1 _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10532__I _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _02739_ _02740_ _02741_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09723_ _04401_ _04407_ _03703_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06935_ _01848_ _01849_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09654_ _02765_ _01651_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06866_ _01780_ _01731_ _01781_ _01783_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_97_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08180__A1 _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07841__I _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08605_ _01690_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05817_ _00825_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06797_ _01717_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09585_ net199 _01615_ _01492_ _01598_ _04267_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_167_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ _03227_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05748_ _00709_ as2650.regs\[6\]\[6\] _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05679_ _00692_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08467_ _01369_ _03171_ _03177_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06494__A1 _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10290__A2 _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ _02187_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08398_ _03114_ _03115_ _03116_ _03118_ _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07349_ net268 _02166_ _02188_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08235__A2 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09432__A1 net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ _03573_ _04934_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output277_I net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09019_ _03706_ _02603_ _03708_ _03710_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_130_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10291_ _04712_ _04867_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09735__A2 _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07237__B _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_126_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09499__A1 _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07751__I _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08171__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11745_ _00529_ clknet_leaf_115_wb_clk_i as2650.stack\[0\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09671__A1 _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09671__B2 _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09678__I _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06485__A1 _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11676_ _00460_ clknet_leaf_17_wb_clk_i as2650.stack\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10627_ _05104_ _05135_ _05137_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09974__A2 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10558_ as2650.stack\[15\]\[6\] _05086_ _05091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06788__A2 _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_126_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10489_ _05016_ _04665_ _04522_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_20_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06830__I _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09726__A2 _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06720_ _01638_ _01645_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08162__A1 _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06651_ as2650.chirp_ptr\[1\] _01586_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_133_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05602_ as2650.indirect_target\[4\] _00599_ _00615_ as2650.PC\[4\] _00616_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_59_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06582_ _01530_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06277__I as2650.cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04046_ _04055_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_133_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ _03043_ _03044_ _03028_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08252_ _02968_ _02983_ _02984_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_1788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07203_ _02058_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ as2650.instruction_args_latch\[14\] _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07134_ net97 net131 _02015_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_65_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09965__A2 _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07976__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06779__A2 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07065_ _01969_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput220 net220 la_data_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput231 net231 last_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10980__B1 _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput242 net242 requested_addr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06016_ _00721_ net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput253 net253 requested_addr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput264 net264 rom_bus_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput275 net275 wbs_dat_o[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput286 net286 wbs_dat_o[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput297 net297 wbs_dat_o[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input36_I io_in[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07967_ _01122_ _01123_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09706_ _04382_ _04385_ _04386_ _04391_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_74_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06918_ _01825_ _01833_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_138_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07898_ _01333_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09637_ as2650.debug_psu\[4\] _02578_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06849_ _00895_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07900__A1 _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06703__A2 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06187__I _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09568_ _01026_ _01656_ net215 _01388_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08519_ _01452_ _03223_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09653__A1 _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09499_ _01129_ _03587_ _01511_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_65_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09653__B2 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11530_ _00314_ clknet_leaf_151_wb_clk_i as2650.stack\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_83_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11461_ _00245_ clknet_leaf_44_wb_clk_i as2650.PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09405__A1 _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06219__A1 _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10412_ _04726_ _04984_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_104_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11392_ _00007_ clknet_leaf_65_wb_clk_i as2650.cycle\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08759__A3 _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07967__A1 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10343_ _04910_ _04861_ _04915_ _04916_ _04917_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_60_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09708__A2 _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_72_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10274_ _04358_ _04796_ _04734_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_72_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08778__S _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_92_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09644__A1 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07430__B _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11728_ _00512_ clknet_leaf_76_wb_clk_i as2650.regs\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_61_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11659_ _00443_ clknet_leaf_78_wb_clk_i as2650.regs\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06473__A4 _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10006__A2 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07958__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08080__B1 as2650.indirect_target\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ as2650.stack\[3\]\[12\] _03495_ _02541_ as2650.stack\[2\]\[12\] _03563_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_55_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07821_ _01429_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_36_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07752_ _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08135__A1 as2650.instruction_args_latch\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06703_ _01605_ net210 _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07683_ _01060_ _01552_ _02451_ _02456_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06697__A1 _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09422_ _04090_ _04091_ _04107_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_75_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06634_ _00697_ net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_94_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09353_ _04035_ _04038_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06565_ as2650.ext_io_addr\[7\] _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09635__A1 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08436__B _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08304_ as2650.instruction_args_latch\[12\] _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_168_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06496_ _01088_ _01458_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09284_ _03966_ _03956_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07110__A2 _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09111__I _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08235_ _02969_ _02620_ _02952_ net198 _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05672__A2 _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08166_ as2650.ivectors_base\[11\] _02852_ _01548_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07117_ net104 net71 _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_82_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08097_ as2650.indirect_target\[9\] _01255_ _02848_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07048_ as2650.stack\[12\]\[14\] _01941_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_164_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__B1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10181__A1 _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08999_ _02787_ _01214_ _03593_ _03596_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__07515__B _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08126__A1 as2650.ivectors_base\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_117_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_117_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_39_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10961_ _05255_ _05267_ _05341_ _05395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_168_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10484__A2 _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10892_ _05301_ _05318_ _05319_ _05331_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_65_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07101__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11513_ _00297_ clknet_leaf_52_wb_clk_i net140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10167__I _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11444_ _00228_ clknet_leaf_37_wb_clk_i as2650.ivectors_base\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11375_ _00171_ clknet_leaf_62_wb_clk_i as2650.insin\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold44_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10326_ _04390_ _04846_ _04900_ _04901_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_123_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10257_ _04723_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10188_ _04725_ _04726_ _04762_ _04766_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__10172__A1 _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07425__B _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__I2 net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06679__A1 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06350_ _01314_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06281_ _00999_ _01039_ net351 _01073_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_44_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08020_ _02770_ _02647_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09087__B _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06603__A1 _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__I as2650.cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09971_ _04597_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08922_ _03588_ _01642_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08356__A1 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08853_ _03543_ _03544_ _03545_ _03546_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_97_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07804_ _02572_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10540__I _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08784_ _03278_ _03479_ _03480_ _03194_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05996_ _00972_ _00979_ _00991_ _00996_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_07735_ _02503_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_139_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08659__A2 _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07666_ net400 _02340_ _02434_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09405_ _03910_ _03926_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06617_ wb_debug_cc _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_14_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07597_ _02373_ _02388_ _02389_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08166__B _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_153_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09336_ _04011_ _04021_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_75_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06548_ _01502_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_35_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09267_ _03945_ _03948_ _03952_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_106_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06479_ _01426_ _01433_ _01435_ _01441_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_4
XANTENNA__08831__A2 _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08218_ _01040_ _02955_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_112_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09198_ _03878_ _03882_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08149_ _00634_ _01440_ _02896_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_1710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07398__A2 _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11160_ as2650.stack\[13\]\[8\] _05536_ _05537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10111_ _04661_ _04687_ _04691_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06070__A2 _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11091_ _05179_ _05487_ _05488_ _05492_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08347__A1 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10042_ _01882_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold30 _02366_ net374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08898__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold41 net463 net385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10450__I _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold52 net76 net396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold63 _00126_ net407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold74 net464 net418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09016__I _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold85 wbs_dat_i[7] net431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold96 wbs_dat_i[9] net442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10944_ as2650.chirpchar\[6\] _05271_ _05379_ _05272_ _05380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_129_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10875_ _04726_ _05315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06375__I _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A2 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_14_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_14_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_152_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05636__A2 _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_97_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11427_ _00211_ clknet_leaf_52_wb_clk_i as2650.instruction_args_latch\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__10625__I _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11358_ _00154_ clknet_leaf_103_wb_clk_i wb_counter\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10309_ _01401_ _01504_ _04734_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_103_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11289_ _00085_ clknet_leaf_1_wb_clk_i net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08889__A2 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05850_ as2650.instruction_args_latch\[0\] _00742_ _00659_ _00857_ _00858_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05781_ _00791_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_99_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07520_ wb_counter\[0\] wb_counter\[1\] wb_counter\[2\] _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08765__I _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07313__A2 _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07451_ _02251_ _02274_ _02276_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11191__I _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06402_ _01366_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05875__A2 _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06285__I _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07382_ _02187_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_146_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09066__A2 _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _01295_ _03807_ _03809_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_161_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06333_ _01299_ _01301_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08274__B1 _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08813__A2 _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09596__I _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09052_ _01343_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06264_ as2650.warmup\[0\] as2650.warmup\[1\] net355 _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_72_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08003_ _02632_ _02759_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10535__I _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06195_ _01163_ _01167_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10384__A1 _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09954_ _00980_ net237 _03105_ _01618_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_146_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07844__I _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08905_ _03594_ _03596_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_5_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10136__A1 _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09885_ as2650.stack\[5\]\[11\] _04540_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08836_ _01905_ _02464_ _03241_ _03530_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_20_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08767_ _02504_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_159_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05979_ _00947_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09829__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07718_ _01873_ _01886_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08698_ _02674_ _03395_ _03397_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_68_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08501__A1 _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07649_ _02423_ _02430_ _02431_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10660_ as2650.regs\[1\]\[6\] _05161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_165_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09319_ _04002_ _04003_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10591_ _05016_ _01970_ _04523_ _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_118_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06815__A1 _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06923__I _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_135_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10445__I _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11212_ _05550_ _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_131_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11143_ _05443_ _05522_ _05526_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_132_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_132_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_133_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11074_ as2650.regs\[7\]\[0\] _05483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10025_ _01800_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08740__B2 as2650.stack\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09296__A2 _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10927_ _05361_ _05362_ _05363_ _05364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10858_ _05296_ _05297_ _05298_ _00871_ _05299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09048__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10789_ as2650.stack\[6\]\[6\] _05238_ _05241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06833__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_1646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06951_ _01864_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10118__A1 _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05793__A1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05902_ as2650.regs\[3\]\[4\] _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09670_ _02676_ _01372_ _03741_ _02658_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06882_ _01784_ _01799_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_141_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08621_ _01792_ _03195_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05833_ as2650.regs\[3\]\[0\] _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_136_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_308 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08552_ _02518_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08495__I _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_319 irq[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_05764_ _00766_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09287__A2 _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07503_ net165 _02305_ _02314_ _02236_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_114_1731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08483_ _02659_ _03187_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05695_ _00708_ _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07434_ net119 _02245_ _02193_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10841__A2 _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07365_ _02174_ _02200_ _02202_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09104_ _03709_ _02615_ _02567_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08798__B2 as2650.stack\[13\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06316_ _01286_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06743__I _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07296_ wb_reset_override _02141_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10265__I _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09035_ _01193_ _01215_ _03726_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_143_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06247_ _01131_ _01219_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input66_I wb_rst_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06178_ _01150_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_106_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09937_ _02739_ _04570_ _04577_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11096__I _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09868_ _04527_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08722__A1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08819_ _03245_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09799_ _01683_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_139_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05822__I _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11761_ _00540_ clknet_leaf_19_wb_clk_i as2650.stack\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10712_ _05078_ _05189_ _05193_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11692_ _00476_ clknet_leaf_79_wb_clk_i as2650.regs\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ _04571_ _05144_ _05148_ _05150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_9_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07749__I _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08789__A1 _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10574_ _01927_ _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_94_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10596__A1 as2650.stack\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__A2 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer8 _00907_ net352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10348__A1 _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10899__A2 _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11126_ _05496_ _05515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_34_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11057_ _05440_ _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10008_ as2650.stack\[4\]\[15\] _04616_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06828__I _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05732__I _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07819__A3 _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__A2 _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06563__I _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07150_ net73 net123 _02025_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06101_ _01077_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10085__I _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07081_ as2650.stack\[11\]\[4\] _01981_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06255__A2 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06032_ _01020_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_105_1708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10339__A1 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08711__C _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_143_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07755__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07983_ _02711_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09722_ _02583_ _04405_ _04406_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06934_ _01786_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09653_ _02765_ _01651_ _01660_ _02769_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06865_ _01782_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08439__B _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08180__A2 _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ as2650.stack\[12\]\[2\] _03305_ _03306_ as2650.stack\[13\]\[2\] _03307_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05816_ _00824_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09584_ as2650.debug_psl\[1\] _04253_ _04265_ _04268_ _04269_ _04270_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_06796_ _01711_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_132_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_121_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08535_ _03195_ _03238_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11067__A2 _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05747_ as2650.regs\[2\]\[6\] _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10814__A2 _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08466_ as2650.ivectors_base\[6\] _03172_ _03175_ _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05678_ _00691_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_161_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09680__A2 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07417_ _02244_ wb_counter\[20\] _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07691__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06494__A2 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08397_ as2650.stack\[15\]\[14\] _02539_ _02542_ as2650.stack\[14\]\[14\] _03117_
+ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_135_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07348_ _02187_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09432__A2 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06246__A2 _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07279_ _02114_ wb_counter\[3\] _02126_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09018_ _03709_ _02602_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output172_I net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ _01626_ _04864_ _04866_ _04719_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_131_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07518__B _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_70_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09499__A2 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_83_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09024__I _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11058__A2 _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09120__A1 _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11744_ _00528_ clknet_leaf_115_wb_clk_i as2650.stack\[0\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10805__A2 _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09671__A2 _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07682__A1 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06485__A2 _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11675_ _00459_ clknet_leaf_18_wb_clk_i as2650.stack\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06383__I _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ as2650.stack\[7\]\[12\] _05136_ _05137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07434__A1 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08631__B1 _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _01852_ _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07985__A2 _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10488_ _04663_ _05038_ _05043_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05748__A1 _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11109_ as2650.stack\[14\]\[5\] _05503_ _05505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06650_ as2650.chirp_ptr\[0\] _01580_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06173__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05601_ _00614_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06581_ _01000_ _01529_ _01273_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08320_ _03034_ _02927_ _03026_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_133_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08251_ as2650.instruction_args_latch\[5\] _02978_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07673__A1 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08870__B1 _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _02057_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06293__I _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08182_ _01998_ as2650.indexed_cyc\[1\] _02915_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07133_ _02018_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06228__A2 _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07064_ _01968_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_144_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput210 net210 la_data_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput221 net221 last_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10980__A1 _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput232 net232 last_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06015_ _01011_ net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput243 net243 requested_addr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10543__I _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput254 net254 requested_addr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput265 net265 wbs_ack_o vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08925__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput276 net276 wbs_dat_o[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_166_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08013__I _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput287 net287 wbs_dat_o[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05739__A1 _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07966_ _02634_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_162_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09705_ _04387_ _04388_ _04389_ _04390_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA_input29_I bus_in_timers[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ _01787_ _01830_ _01832_ _01798_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_74_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07897_ _02658_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08153__A2 _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09350__A1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09636_ _01559_ _02465_ _04321_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_39_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06848_ _00610_ _01741_ _01766_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__06164__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09567_ _01855_ _03744_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05911__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06779_ _01509_ _01699_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09102__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ _00594_ _01473_ _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09498_ _04156_ _04182_ _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_136_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09653__A2 _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__I _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ as2650.ivectors_base\[0\] _03165_ _02809_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11460_ _00244_ clknet_leaf_42_wb_clk_i as2650.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_22_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10411_ _04389_ _04846_ _04982_ _04983_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_116_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11391_ _00006_ clknet_leaf_68_wb_clk_i as2650.cycle\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_145_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_76_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07967__A2 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10342_ _01461_ _01505_ _04710_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_60_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10273_ _04736_ _04737_ _01410_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_72_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05993__A4 _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_39_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_39_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10402__B _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06378__I _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08593__I _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09644__A2 _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06458__A2 _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11727_ _00511_ clknet_4_15__leaf_wb_clk_i as2650.regs\[0\]\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_100_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11658_ _00442_ clknet_leaf_95_wb_clk_i as2650.regs\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07002__I _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10609_ _05088_ _05123_ _05126_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08604__B1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11589_ _00373_ clknet_leaf_8_wb_clk_i as2650.stack\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08080__A1 as2650.instruction_args_latch\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05969__A1 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08080__B2 _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10962__A1 _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08907__A1 _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10714__A1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09580__A1 _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ _01315_ _02588_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_104_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07672__I _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06394__A1 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11355__CLK clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ _02519_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06702_ net241 _01602_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08135__A2 _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ net230 _02452_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07194__I0 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09421_ _03915_ _04106_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06633_ _00787_ net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09352_ _04036_ _04037_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06564_ as2650.io_bus_we _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_48_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08303_ _02933_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06449__A2 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09283_ _03929_ _03936_ _03968_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06495_ _01247_ _01451_ _01454_ _01457_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_16_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07110__A3 _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08234_ _01251_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08165_ as2650.indirect_target\[15\] _02909_ _02910_ _02723_ _02630_ _02911_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_126_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07116_ _01999_ _02002_ _02004_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08071__A1 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08096_ _01723_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10953__A1 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07047_ _01953_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09571__A1 _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__B2 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08998_ _03685_ _03687_ _03689_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10181__A2 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output135_I net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07949_ _01468_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10222__B _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10960_ _05261_ _05391_ _05392_ _05394_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07185__I0 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09619_ _04293_ _04302_ _04303_ _04304_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_104_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10891_ _05301_ _05330_ _05331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_65_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_157_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_157_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07637__A1 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10448__I _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08834__B1 _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11512_ _00296_ clknet_leaf_66_wb_clk_i net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_136_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11443_ _00227_ clknet_leaf_37_wb_clk_i as2650.ivectors_base\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06860__A2 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08062__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11374_ _00170_ clknet_leaf_62_wb_clk_i as2650.insin\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10325_ _02731_ _04898_ _04845_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold37_I net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10256_ _04832_ _04833_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_101_1722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09562__A1 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06376__A1 _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10187_ _04763_ _04765_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10172__A2 _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_89_wb_clk_i_I clknet_4_10__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07176__I0 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06679__A2 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07441__B _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05740__I _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09617__A2 _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06280_ _01251_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06300__A1 _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08053__A1 as2650.indirect_target\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09087__C _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06064__B1 _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09970_ _04594_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_122_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08921_ _03611_ _03612_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_21_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08356__A2 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ as2650.stack\[15\]\[11\] _01692_ _01968_ as2650.stack\[14\]\[11\] _02520_
+ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_100_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07803_ _01254_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08783_ _01878_ _03195_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05995_ net236 _00987_ _00993_ _00995_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_93_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07734_ _02502_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07167__I0 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11112__A1 _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07665_ wb_counter\[30\] _02443_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09404_ _03912_ _03925_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_157_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06616_ _01559_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_157_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07596_ net386 _02376_ _02385_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09608__A2 as2650.debug_psu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09335_ _01015_ _01495_ _01489_ net190 _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_146_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06547_ _00969_ _00998_ _01075_ _01081_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_36_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09084__A3 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09266_ _03949_ _03950_ _03951_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06478_ _01434_ _01431_ _01439_ _01440_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_47_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08217_ _02954_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06842__A2 _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09197_ _03882_ _03878_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__07577__I _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _02895_ _01440_ _02660_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08079_ _02708_ _01456_ _02831_ _02724_ as2650.indirect_target\[8\] _02832_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__09792__B2 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10110_ as2650.stack\[3\]\[14\] _04688_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output252_I net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06070__A3 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11090_ as2650.regs\[7\]\[7\] _05492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10041_ _04643_ _04636_ _04644_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold20 _00125_ net364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold31 _00139_ net375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold42 net79 net386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold53 net448 net397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold64 net436 net408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold75 net446 net419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold86 wbs_dat_i[3] net432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold97 wbs_dat_i[28] net443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05581__A2 as2650.cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07858__A1 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10943_ _05377_ _05378_ _05304_ _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10874_ _05295_ _05299_ _05300_ _05314_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_109_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08807__B1 _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11426_ _00210_ clknet_leaf_65_wb_clk_i as2650.instruction_args_latch\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06391__I net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_54_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09783__A1 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11357_ _00153_ clknet_leaf_101_wb_clk_i wb_counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10308_ _04736_ _04883_ _01404_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11288_ _00084_ clknet_leaf_1_wb_clk_i net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_52_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08338__A2 _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _02922_ _04753_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07436__B _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06340__B _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05780_ _00790_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_76_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08510__A2 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07450_ net283 _02256_ _02275_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06401_ _01280_ _01365_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07381_ _02211_ wb_counter\[15\] _02216_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05875__A3 _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09877__I _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09120_ _01780_ _02739_ _03808_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06332_ _00647_ _01300_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_127_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09051_ _01204_ _01214_ _01398_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__10081__A1 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06263_ _01088_ _01235_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08002_ _02756_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06380__S0 _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08026__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06194_ _01166_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_83_1743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06588__A1 _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09953_ _01603_ _04587_ _03051_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_99_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10551__I _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08904_ _01667_ _03587_ _03595_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_146_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09884_ _01913_ _04539_ _04543_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07001__A2 _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08835_ _01909_ _03375_ _03529_ _03242_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_100_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ as2650.stack\[3\]\[8\] _03461_ _03462_ as2650.stack\[2\]\[8\] _03463_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_159_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05978_ net236 _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_input11_I bus_in_serial_ports[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07717_ as2650.stack\[3\]\[13\] _01693_ _01969_ as2650.stack\[2\]\[13\] _02486_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_101_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08697_ _03090_ _03396_ _02667_ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08177__B _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07648_ net90 _02426_ _02418_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06512__A1 _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07579_ wb_counter\[13\] _02374_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_3_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09318_ _04002_ _04003_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08265__A1 as2650.instruction_args_latch\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10590_ _05112_ _05105_ _05113_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_149_Left_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08624__C _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09249_ _00766_ _01016_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07100__I _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11211_ _05548_ _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_131_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09765__A1 _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11142_ as2650.stack\[13\]\[1\] _05524_ _05526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11073_ _05481_ _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_158_Left_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10024_ _04631_ _04625_ _04632_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08740__A2 _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06751__A1 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__I _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_101_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_101_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10926_ as2650.chirpchar\[5\] _05267_ _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10857_ _05285_ _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_45_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10850__A3 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_167_Left_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_99_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08256__A1 as2650.instruction_args_latch\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10788_ _05088_ _05237_ _05240_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08008__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08559__A2 _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11409_ _00193_ clknet_leaf_48_wb_clk_i as2650.indirect_target\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06950_ _01862_ _01863_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10118__A2 _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I bus_in_gpios[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05901_ _00841_ _00906_ _00829_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06881_ _01787_ _01792_ _01794_ _01798_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_141_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08620_ _03085_ _03321_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05832_ _00829_ _00840_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06742__A1 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ as2650.stack\[7\]\[1\] _03244_ _03254_ as2650.stack\[6\]\[1\] _03255_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_309 io_oeb[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_05763_ _00758_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_37_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07502_ net100 _02058_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08482_ net204 _03067_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05694_ _00707_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07433_ _02251_ _02260_ _02261_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07364_ _02201_ _02141_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09103_ _01772_ _02944_ _03791_ _03792_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_45_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06315_ _01131_ _01276_ _01216_ _01285_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_116_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10546__I _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07295_ net69 _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _01195_ _02563_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_14_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06246_ _01184_ _01202_ _01218_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_5_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09747__A1 _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06177_ _01148_ _01149_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_148_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07855__I _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input59_I rom_bus_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10281__I _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ net143 _04576_ _04572_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10109__A2 _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09867_ _04525_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08722__A2 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _01917_ _03512_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07590__I _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09798_ _04429_ _04478_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output215_I net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _03107_ _02819_ _03399_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11760_ _00539_ clknet_leaf_99_wb_clk_i as2650.regs\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08486__A1 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10711_ as2650.stack\[8\]\[1\] _05191_ _05193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11691_ _00475_ clknet_leaf_95_wb_clk_i as2650.regs\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_137_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08238__A1 as2650.instruction_args_latch\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10642_ _05148_ _05149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _05100_ _05095_ _05101_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer9 _00906_ net353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_wire299_I net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06264__A3 net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11125_ _05494_ _05514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08961__A2 _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09980__I _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11056_ _05438_ _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10007_ _01954_ _04615_ _04619_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06724__A1 net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07005__I as2650.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10909_ as2650.regs\[4\]\[3\] _05335_ _05347_ _05301_ _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_39_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09977__A1 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10366__I _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06100_ _01076_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10587__A2 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07080_ _01974_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06031_ _01019_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09729__A1 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07675__I _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09095__C _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08952__A2 _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07982_ _02660_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06963__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05766__A2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06933_ _01844_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09721_ _02583_ _04400_ _04354_ _02586_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_138_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _02769_ _01660_ _04335_ _04337_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_59_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06864_ _01711_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08603_ _03250_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05815_ _00823_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09583_ as2650.debug_psl\[1\] _04266_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06795_ _01715_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08534_ _03237_ _01744_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05746_ _00757_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08468__A1 as2650.ivectors_base\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__B2 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08465_ _01351_ _03171_ _03176_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05677_ _00690_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_148_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07416_ _02192_ _01924_ _02246_ _02170_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_50_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06494__A3 _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08396_ _02519_ _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_169_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__A1 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07347_ _02073_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10276__I _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07278_ _02116_ _02123_ _02125_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_147_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09017_ _02590_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06229_ _01189_ _01201_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_83_1370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output165_I net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06954__A1 _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10750__A2 _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09919_ _04562_ _01657_ _04566_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_70_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06929__I as2650.PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_83_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09120__A2 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11743_ _00527_ clknet_leaf_116_wb_clk_i as2650.stack\[0\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11674_ _00458_ clknet_leaf_21_wb_clk_i as2650.stack\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09959__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10625_ _05117_ _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_148_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07434__A2 _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold67_I _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10556_ _05088_ _05085_ _05089_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10487_ as2650.stack\[2\]\[15\] _05039_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08395__B1 _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06945__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10741__A2 _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ _05449_ _05502_ _05504_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11039_ as2650.stack\[0\]\[7\] _05451_ _05458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08698__A1 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05600_ _00593_ _00595_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_34_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06580_ _01528_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05920__A2 _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08250_ _02969_ _02577_ _02976_ net201 _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07673__A2 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07201_ _02056_ _02008_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05684__A1 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ _02916_ _02923_ _02925_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_9_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_70_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07132_ net94 net130 _02015_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07063_ _01967_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput200 net200 la_data_out[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06523__B _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput211 net211 la_data_out[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05918__I _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput222 net222 last_addr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06014_ _00988_ _00974_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput233 net233 last_addr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_144_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput244 net244 requested_addr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_122_1820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput255 net255 requested_addr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_151_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput266 net266 wbs_dat_o[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput277 net277 wbs_dat_o[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_166_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput288 net288 wbs_dat_o[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09834__B _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06936__A1 _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07965_ _01305_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_96_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09704_ net4 net12 net28 net20 _04383_ _01520_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_06916_ _01831_ _01793_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07896_ _02645_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08689__B2 _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09125__I _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08169__C _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _01950_ _01577_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06847_ _01742_ _01765_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06778_ _01698_ _01284_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_91_1661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09566_ _03160_ _03768_ _03725_ _04197_ _04251_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_151_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09102__A2 _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05729_ _00588_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08517_ _03217_ _03221_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07113__A1 _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09497_ _01229_ _01285_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_108_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08448_ _03163_ _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_81_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08379_ _01257_ _02934_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_22_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10410_ _02790_ _04898_ _04845_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11390_ _00016_ clknet_leaf_65_wb_clk_i as2650.cycle\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07416__A2 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output282_I net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09728__C _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10341_ _04360_ _04793_ _04811_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06624__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10272_ _04803_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_72_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08916__A2 _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_79_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_1578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10239__A1 _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08807__C _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11726_ _00510_ clknet_leaf_81_wb_clk_i as2650.regs\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08852__B2 as2650.stack\[14\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11657_ _00441_ clknet_leaf_93_wb_clk_i as2650.regs\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10608_ as2650.stack\[7\]\[5\] _05124_ _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11588_ _00372_ clknet_leaf_11_wb_clk_i as2650.stack\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10411__A1 _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08080__A2 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10539_ _05071_ _05074_ _05077_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05969__A2 net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10962__A2 _05395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08907__A2 _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06918__A1 _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07953__I _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10714__A2 _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09580__A2 _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09707__I1 net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07750_ _02518_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_75_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06701_ _01550_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07681_ _02454_ _02455_ _02004_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07194__I1 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09420_ _04093_ _04105_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06632_ _00814_ net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_152_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06563_ _01516_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09351_ net220 _01490_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09096__A1 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06518__B _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08302_ _03025_ _03027_ _03028_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09282_ net217 net220 _03934_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06494_ _01089_ _01322_ _01456_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08843__A1 _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08233_ _02572_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10650__A1 _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10650__B2 _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08164_ _01335_ _02843_ _00644_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_145_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07115_ _02003_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10402__A1 _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10554__I _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08095_ _02846_ _02740_ _02741_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_113_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__B _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07046_ _01949_ _01843_ _01952_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_110_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_164_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06909__A1 _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07863__I _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input41_I io_in[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08997_ _03653_ _03688_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _02001_ _02706_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09323__A2 _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07879_ _02639_ _02640_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_output128_I net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07185__I1 net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09618_ _01559_ _02943_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10890_ _05328_ _05329_ _05330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_104_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05896__A1 _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09549_ _04232_ _03826_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09087__A1 _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11511_ _00295_ clknet_leaf_69_wb_clk_i net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_53_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10641__A1 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09739__B _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_152_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_126_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_126_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11442_ _00226_ clknet_leaf_37_wb_clk_i as2650.ivectors_base\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06942__I _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11373_ _00169_ clknet_leaf_30_wb_clk_i as2650.debug_psu\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10324_ _04882_ _04894_ _04897_ _04899_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_132_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10255_ _04247_ _04831_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__07773__I _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09562__A2 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10186_ _04387_ _04764_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06376__A2 _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08770__B1 _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06389__I _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07176__I1 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09078__A1 _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07441__C _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11709_ _00493_ clknet_leaf_22_wb_clk_i as2650.stack\[6\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06852__I as2650.debug_psl\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11188__A2 _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06064__B2 as2650.cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__A2 _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08920_ _01124_ _03585_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10699__A1 _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ as2650.stack\[12\]\[11\] _03137_ _03138_ as2650.stack\[13\]\[11\] _03545_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11472__CLK clknet_4_12__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07802_ _02483_ _02558_ _02570_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_100_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05994_ net225 _00961_ _00994_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
Xclkbuf_1_1__f__01549_ clknet_0__01549_ clknet_1_1__leaf__01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08782_ _03374_ _03457_ _03478_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07733_ _02501_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_139_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07167__I1 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ wb_counter\[29\] _02440_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09403_ _03981_ _04082_ _04087_ _04088_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_157_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06615_ as2650.debug_psl\[6\] _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07595_ wb_counter\[16\] _02387_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10549__I _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09069__A1 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09608__A3 net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06546_ wb_io3_test net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_09334_ _04018_ _04019_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08816__A1 _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08816__B2 _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10623__A1 _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06477_ _01300_ _01424_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_8_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09265_ _03871_ _00825_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08216_ _01336_ _01332_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _03879_ _03880_ _03881_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_47_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10284__I _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ _02894_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08044__A2 _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09241__A1 _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08078_ _02794_ _02830_ _02804_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07029_ _01849_ _01936_ _01937_ _01842_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_12_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10040_ as2650.stack\[10\]\[7\] _04637_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output245_I net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__A2 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold21 net432 net365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_95_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold32 net440 net376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold43 net441 net387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold54 net77 net398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold65 _02028_ net409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold76 net461 net420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold87 _02334_ net433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07307__A1 net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold98 wbs_adr_i[22] net444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_93_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08504__B1 _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11103__A2 _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05581__A3 as2650.cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10942_ net193 _04772_ _05378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10459__I _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10873_ _05301_ _05313_ _05314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08807__A1 _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11425_ _00209_ clknet_leaf_66_wb_clk_i as2650.instruction_args_latch\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11356_ _00152_ clknet_leaf_101_wb_clk_i wb_counter\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09783__A2 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07794__A1 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10307_ _04703_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11287_ _00083_ clknet_leaf_1_wb_clk_i net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_52_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_94_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_94_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_123_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10238_ _01415_ _04792_ _04812_ _04813_ _04815_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_TAPCELL_ROW_52_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07546__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_23_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_23_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10169_ _04746_ _04747_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06400_ _01180_ _01364_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_119_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07380_ _02212_ _02214_ _02215_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09846__I0 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06331_ _01209_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_70_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09050_ _01193_ _01215_ _03726_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06262_ _01089_ _01094_ _01234_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold119_I wbs_dat_i[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ as2650.indirect_target\[4\] _02757_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06380__S1 _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06193_ _01142_ _01165_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_108_1729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06588__A2 _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09952_ net235 _04586_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08903_ _03589_ _01669_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ as2650.stack\[5\]\[10\] _04540_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_10__f_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08734__B1 _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08834_ _03337_ _03513_ _03528_ _03324_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08765_ _03245_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05977_ net223 net242 _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_169_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_159_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07716_ _02484_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_101_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _03073_ _03087_ _03089_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_101_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10844__A1 _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07647_ wb_counter\[26\] _02429_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_152_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ wb_counter\[11\] wb_counter\[12\] _02364_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_113_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09317_ _03937_ _03954_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_36_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06529_ _00856_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__A1 _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09248_ _03930_ _03932_ _03933_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output195_I net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09179_ _03702_ _03865_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11210_ _05467_ _05562_ _05567_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11141_ _05436_ _05522_ _05525_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05836__I _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08212__I _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11072_ _05168_ _05479_ _05481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07528__A1 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput100 net389 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10023_ as2650.stack\[10\]\[2\] _04627_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07272__B net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10925_ net192 _04933_ _05271_ _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_141_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_141_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold97_I wbs_dat_i[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10856_ _05284_ _05297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10787_ as2650.stack\[6\]\[5\] _05238_ _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_41_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10063__A2 _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11408_ _00192_ clknet_leaf_46_wb_clk_i as2650.indirect_target\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11339_ _00135_ clknet_leaf_143_wb_clk_i wb_counter\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05900_ _00883_ _00905_ _00900_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_118_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06880_ _01797_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_141_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08192__A1 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05831_ _00661_ _00834_ _00839_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06577__I _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08550_ _03245_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05762_ _00680_ _00771_ _00772_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_76_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10320__C _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07501_ _02312_ net363 _02309_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10826__A1 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08481_ _02640_ net204 _03067_ _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05693_ _00691_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09692__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09888__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07432_ net280 _02256_ _02249_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07363_ _01808_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06526__B _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09102_ _01769_ _03747_ _02944_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06314_ _01167_ _01284_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_31_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07294_ net133 _02139_ _02122_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06245_ _01208_ _01216_ _01217_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_5_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09033_ _03724_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11003__A1 _05384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06176_ as2650.insin\[6\] _01095_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09747__A2 _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09128__I _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09935_ _01464_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08032__I _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09866_ _01801_ _04526_ _04532_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08817_ _01877_ _01890_ _03459_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09797_ _01683_ _04476_ _04477_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07930__A1 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07930__B2 _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06487__I _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08748_ _03237_ _01865_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_124_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output110_I net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10817__A1 _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08486__A2 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output208_I net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ as2650.stack\[4\]\[5\] _02491_ _02498_ as2650.stack\[5\]\[5\] _03204_ _03379_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_95_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06497__A1 _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10710_ _05071_ _05189_ _05192_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11690_ _00474_ clknet_leaf_87_wb_clk_i as2650.chirpchar\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_81_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10737__I _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10641_ _01808_ _05147_ _05148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_137_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10572_ as2650.stack\[15\]\[10\] _05096_ _05101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_165_Right_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07111__I _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07997__A1 _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06421__A1 _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11124_ _05467_ _05508_ _05513_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11055_ _01939_ _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_34_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__I _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10006_ as2650.stack\[4\]\[14\] _04616_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09910__A2 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A1 _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06488__A1 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06488__B2 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _05345_ _05346_ _05347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09426__A1 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10839_ _05278_ _05279_ _05280_ _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_17_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09977__A2 _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07021__I _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__B2 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07956__I _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06030_ _00846_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09729__A2 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06412__A1 _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07981_ _02731_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_10_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_26_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09720_ _01564_ _02991_ _03718_ _04404_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06932_ _01742_ _01846_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08165__A1 as2650.indirect_target\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08165__B2 _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _04334_ _04336_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06863_ net214 _01732_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06715__A2 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07912__A1 _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08602_ _03248_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05814_ _00789_ as2650.regs\[4\]\[3\] _00822_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_09582_ _04253_ _04267_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06794_ _01714_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_116_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08533_ _03229_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05745_ _00756_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09665__A1 _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06479__A1 _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08464_ as2650.ivectors_base\[5\] _03172_ _03175_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05676_ _00689_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ net116 _02245_ _02193_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10557__I _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08395_ as2650.stack\[12\]\[14\] _02534_ _02537_ as2650.stack\[13\]\[14\] _03116_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_169_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07346_ _02181_ wb_counter\[11\] _02185_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07277_ web_behavior\[1\] _02124_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09016_ _03707_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06228_ _01194_ _01200_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_131_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06159_ _01119_ _01105_ _01106_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_79_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _04563_ net152 _04564_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_4_13__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09849_ _04520_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_87_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06706__A2 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_83_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11742_ _00526_ clknet_leaf_136_wb_clk_i as2650.stack\[0\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11673_ _00457_ clknet_leaf_100_wb_clk_i as2650.regs\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09408__A1 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10624_ _05115_ _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10555_ as2650.stack\[15\]\[5\] _05086_ _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08631__A2 _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10486_ _04661_ _05038_ _05042_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09991__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11107_ as2650.stack\[14\]\[4\] _05503_ _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07217__S _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11038_ _01868_ _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07370__A2 _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__A1 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08870__A2 _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ net69 _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11206__A1 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05684__A2 _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08180_ _01241_ _02924_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07131_ _02017_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06590__I _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold101_I wbs_dat_i[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07062_ _01966_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_109_1643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput201 net201 la_data_out[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06013_ _01010_ net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06523__C _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput212 net212 la_data_out[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_103_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput223 net223 last_addr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput234 net234 last_addr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput245 net245 requested_addr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput256 net355 reset_out vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_34_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput267 net267 wbs_dat_o[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput278 net278 wbs_dat_o[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput289 net289 wbs_dat_o[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07964_ _02710_ _02719_ _02721_ _02722_ _01526_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_96_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08138__A1 as2650.ivectors_base\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09703_ net7 net15 net31 net23 _04383_ _04384_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_06915_ _01826_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07895_ _02656_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09886__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08689__A2 _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09634_ _01558_ _00687_ _04319_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06846_ _01764_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_121_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09565_ _03780_ _03781_ _04210_ _04250_ _03724_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_06777_ _01196_ _01164_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_116_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09638__A1 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_43_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08466__B _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08516_ _01721_ _02482_ _03220_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05728_ _00590_ _00740_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_37_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09496_ _04157_ _04159_ _04181_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_38_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10287__I _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08447_ _03163_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05659_ _00672_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_110_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_142_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08378_ _02895_ _03099_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_119_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07329_ _02147_ _01558_ _02169_ _02170_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08613__A2 _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09810__A1 _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06624__A1 wb_debug_cc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ _04808_ _04913_ _04914_ _04848_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_76_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__C _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_52_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10271_ _04847_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_72_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_128_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07545__B _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08220__I _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10487__A2 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_61_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09629__A1 _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07104__A2 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_48_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_48_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_70_1779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11725_ _00509_ clknet_leaf_76_wb_clk_i as2650.regs\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05666__A2 _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06863__A1 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11656_ _00440_ clknet_leaf_91_wb_clk_i as2650.regs\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_61_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08823__C _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10607_ _05084_ _05123_ _05125_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08604__A2 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11587_ _00371_ clknet_leaf_8_wb_clk_i as2650.stack\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09801__A1 _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10538_ as2650.stack\[15\]\[0\] _05076_ _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_1831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10469_ _05018_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09565__B1 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10175__A1 _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05754__I _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09707__I2 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06700_ _01612_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ net229 _01628_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06631_ _00862_ net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_137_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__B _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09350_ _01496_ _04027_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06585__I _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06562_ _01515_ _01246_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_48_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08301_ _02003_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06518__C _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09281_ _03956_ _03966_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06493_ _01455_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_145_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08232_ _02949_ _02967_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _02689_ _02635_ _02653_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06067__C1 _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07114_ _01086_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08094_ as2650.instruction_args_latch\[9\] _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07045_ _01950_ _01770_ _01951_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_144_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08359__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09020__A2 _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_1369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08996_ _03594_ _03596_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_input34_I io_in[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07947_ _02638_ _02701_ _02704_ _02705_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_58_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06790__B1 _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_108_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07878_ _02602_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09617_ _01429_ _01201_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06829_ _01748_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_1779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_104_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09548_ _04232_ _03634_ _04233_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_65_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09087__A2 _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07098__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09479_ _04008_ _04080_ _04081_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11510_ _00294_ clknet_leaf_68_wb_clk_i net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_117_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06845__A1 _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10641__A2 _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _00225_ clknet_leaf_37_wb_clk_i as2650.ivectors_base\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11372_ _00168_ clknet_leaf_70_wb_clk_i net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10323_ _01404_ _04758_ _04898_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05820__A2 as2650.instruction_args_latch\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10254_ _04827_ _04828_ _04829_ _04831_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__10480__I _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10185_ _04707_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05574__I as2650.cycle\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05584__A1 as2650.relative_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08522__A1 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09078__A2 _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11708_ _00492_ clknet_leaf_22_wb_clk_i as2650.stack\[6\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10632__A2 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08553__C _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11639_ _00423_ clknet_leaf_14_wb_clk_i as2650.stack\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_150_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10396__A1 _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06064__A2 _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07261__A1 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10935__A3 _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09002__A2 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08850_ as2650.stack\[8\]\[11\] _02533_ _02536_ as2650.stack\[9\]\[11\] _03131_ _03544_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07801_ _02569_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08761__A1 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08781_ _01879_ _02464_ _03477_ _01258_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05993_ _00973_ _00983_ _00955_ _00964_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_34_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ as2650.debug_psu\[2\] _01686_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07663_ _02332_ _02441_ _02442_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09402_ _04084_ _04086_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06614_ _01557_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_157_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07594_ wb_counter\[14\] wb_counter\[15\] _02379_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09069__A2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07204__I _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_9_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09333_ _01501_ _01020_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06545_ _01501_ net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08816__A2 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ _01027_ _00815_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06476_ _01438_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08215_ _01252_ _02603_ net195 _02952_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_118_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10565__I _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09195_ _00790_ _00824_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05659__I _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08146_ _02893_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07252__A1 _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08077_ _02826_ _02829_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_144_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__I _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09529__B1 _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07028_ _01934_ _01786_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold22 net97 net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold33 net74 net377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_95_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output238_I net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ _03621_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold44 net75 net388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold55 net456 net399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold66 wbs_adr_i[20] net410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold77 net454 net421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold88 wbs_dat_i[31] net434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold99 wbs_dat_i[6] net445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__07307__A2 _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10941_ _03416_ _05321_ _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06515__B1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10311__A1 _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10872_ _05311_ _04318_ _05312_ _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07114__I _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08807__A2 _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09480__A2 _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11424_ _00208_ clknet_leaf_68_wb_clk_i as2650.instruction_args_latch\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11355_ _00151_ clknet_4_8__leaf_wb_clk_i wb_counter\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold42_I net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10306_ _04757_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_56_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11286_ _00082_ clknet_leaf_150_wb_clk_i net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_123_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10237_ _04814_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_98_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10168_ _04287_ _04744_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10099_ _04649_ _04681_ _04684_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_63_wb_clk_i clknet_4_13__leaf_wb_clk_i clknet_leaf_63_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_156_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10853__A2 _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06330_ as2650.instruction_args_latch\[15\] _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_152_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06261_ _01089_ _01223_ _01233_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_115_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08000_ _02679_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06192_ _01164_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_83_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10369__B2 _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07234__A1 _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09951_ _01544_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_42_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08902_ _02786_ _01227_ _03593_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_21_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09882_ _01899_ _04539_ _04542_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_146_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06103__I _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _03522_ _03527_ _03267_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08764_ _03210_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05976_ _00978_ net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_159_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_159_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07715_ _02472_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11097__A2 _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08695_ _03372_ _03373_ _03394_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_101_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07646_ _02428_ _02424_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_62_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10844__A2 _05258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06512__A3 _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07577_ _02357_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09316_ _03992_ _04000_ _04001_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06528_ _01469_ _01476_ _01487_ _01488_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06773__I _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06276__A2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09247_ _00913_ _00825_ _03931_ _01498_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_88_1656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06459_ _01342_ _01421_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09178_ _03704_ _03864_ _03849_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output188_I net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _02853_ _02867_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_131_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11140_ as2650.stack\[13\]\[0\] _05524_ _05525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_92_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05787__A1 _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10780__A1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11071_ _05479_ _05480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_1730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07109__I _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07528__A2 _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput101 net369 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10022_ _01776_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09752__C _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09150__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10924_ _03386_ _05266_ _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10855_ _04832_ _04833_ _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_45_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10599__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10786_ _05084_ _05237_ _05239_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__A1 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_110_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11407_ _00191_ clknet_leaf_46_wb_clk_i as2650.indirect_target\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08831__C _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08964__A1 _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11338_ _00134_ clknet_leaf_144_wb_clk_i wb_counter\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11269_ _00065_ clknet_leaf_137_wb_clk_i net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__08716__A1 _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08192__A2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05830_ _00811_ as2650.instruction_args_latch\[3\] _00613_ _00838_ _00839_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06858__I _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05761_ _00705_ net202 _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05950__A1 _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07500_ net362 _02307_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08480_ _00722_ _03179_ _03185_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05692_ _00705_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09692__A2 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07431_ _02244_ wb_counter\[22\] _02259_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07362_ net126 _02199_ _02175_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09101_ _03729_ _03769_ _03785_ _03790_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06313_ _01278_ _01283_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07455__A1 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07293_ _02118_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_99_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09032_ _01215_ _03716_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06244_ _01115_ _01209_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_115_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11003__A2 _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06175_ _00664_ _01147_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_148_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09934_ _02716_ _04570_ _04575_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09865_ as2650.stack\[5\]\[3\] _04528_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08816_ _02859_ _03053_ _03510_ _03502_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07373__B _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09796_ _01684_ _03143_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08747_ _01860_ _03283_ _03444_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05959_ _00944_ _00633_ _00962_ _00963_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XANTENNA__05941__A1 _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_124_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09132__A1 _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08678_ as2650.stack\[7\]\[5\] _03200_ _02511_ as2650.stack\[6\]\[5\] _03378_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10817__A2 _05258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06497__A2 _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07629_ wb_counter\[22\] _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10640_ _04693_ _04694_ _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_137_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10571_ _01912_ _05100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09747__C _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_98_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11123_ as2650.stack\[14\]\[11\] _05509_ _05513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09763__B _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11054_ _05467_ _05460_ _05468_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ _01947_ _04615_ _04618_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05582__I _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__B2 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10808__A2 _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08826__C _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07685__A1 _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10907_ _04480_ _02580_ _05280_ _05346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_156_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10838_ _05262_ _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_27_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__A1 net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10769_ _05179_ _05222_ _05223_ _05227_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_82_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08842__B _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08561__C _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09729__A3 _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06362__B _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07980_ _01335_ _02737_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06931_ _01845_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09650_ _02827_ _01669_ _04333_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06862_ _01779_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA__06176__A1 as2650.insin\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08601_ as2650.stack\[8\]\[2\] _03302_ _03303_ as2650.stack\[9\]\[2\] _03294_ _03304_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05813_ _00753_ _00821_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_145_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_1699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09581_ _01667_ _03855_ _04266_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06793_ _01685_ _01694_ _01713_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_91_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08532_ _03186_ _03079_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09114__B2 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05744_ _00755_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08463_ _03174_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08873__B1 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05675_ as2650.debug_psl\[4\] _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07414_ _02117_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ as2650.stack\[8\]\[14\] _02527_ _02530_ as2650.stack\[9\]\[14\] _02506_ _03115_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_clkbuf_leaf_132_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07345_ _02174_ _02182_ _02184_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_11_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07276_ _02056_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_104_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09015_ _01183_ _02565_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_60_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06227_ _01199_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_1384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input64_I rom_bus_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08928__A1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06158_ _01130_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_83_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10735__A1 as2650.stack\[8\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06089_ _01067_ net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09917_ _04562_ _01648_ _04565_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_96_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09848_ net48 as2650.irqs_latch\[6\] _01516_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_126_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07903__A2 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output220_I net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09779_ _04443_ _04450_ _03128_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09105__A1 _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07667__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _00525_ clknet_leaf_130_wb_clk_i as2650.stack\[0\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11672_ _00456_ clknet_leaf_100_wb_clk_i as2650.regs\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07122__I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10623_ _05102_ _05129_ _05134_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_27_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11215__A2 _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08092__A1 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10554_ _01834_ _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10974__A1 _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06642__A2 _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10485_ as2650.stack\[2\]\[14\] _05039_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08919__A1 _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10726__A1 _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_36_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08395__A2 _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11106_ _05496_ _05503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__B _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11650__CLK clknet_leaf_92_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11037_ _05455_ _05450_ _05456_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11151__A1 _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08698__A3 _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08556__C _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07658__A1 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08855__B1 _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07032__I _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07130_ net83 net129 _02015_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08083__A1 as2650.ivectors_base\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__I0 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07061_ _01965_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_152_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06012_ _00976_ _00992_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput202 net202 la_data_out[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_70_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput213 net213 la_data_out[32] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_105_1508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput224 net224 last_addr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_3_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput235 net235 last_addr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput246 net246 requested_addr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_45_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput257 net257 rom_bus_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09583__A1 as2650.debug_psl\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput268 net268 wbs_dat_o[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput279 net279 wbs_dat_o[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_166_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10193__A2 _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07963_ _01450_ as2650.irqs_latch\[6\] as2650.irqs_latch\[7\] _02722_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_09702_ net6 net30 net14 net22 as2650.ext_io_addr\[6\] _01518_ _04388_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_06914_ _01829_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09335__B2 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07894_ _02655_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06111__I _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ _01872_ _00687_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06845_ _00610_ _01763_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_121_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09564_ _04216_ _04249_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06776_ _01696_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09638__A2 _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08515_ _03198_ _03199_ _03219_ _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05727_ _00620_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07649__A1 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10568__I _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ _04160_ _04162_ _04180_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_78_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07113__A3 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08446_ _03162_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05658_ net225 net224 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_147_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08377_ _03030_ _03098_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_34_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05589_ as2650.relative_cyc as2650.indirect_cyc _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_119_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07877__I _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07328_ _02112_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11523__CLK clknet_4_15__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10956__A1 _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06624__A2 _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ wb_counter\[2\] _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_76_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10270_ _01728_ _03730_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_89_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07888__B2 _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11862__I net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06560__A1 _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09629__A2 _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11724_ _00508_ clknet_leaf_81_wb_clk_i as2650.regs\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11655_ _00439_ clknet_leaf_91_wb_clk_i as2650.regs\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_88_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_88_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10606_ as2650.stack\[7\]\[4\] _05124_ _05125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11586_ _00370_ clknet_leaf_9_wb_clk_i as2650.stack\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10537_ _05075_ _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_17_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _04643_ _05026_ _05031_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09565__A1 _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10399_ _03855_ _04971_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08411__I _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11124__A1 _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06630_ _00844_ net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_75_1669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06561_ _01084_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08828__B1 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08300_ _03007_ as2650.instruction_args_latch\[11\] _03026_ _03027_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09280_ _03959_ _03960_ _03965_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_129_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06492_ _01260_ _01268_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08231_ as2650.instruction_args_latch\[2\] _02950_ _02966_ _02958_ _02967_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_144_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06815__B _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07697__I _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08162_ _02899_ _02747_ _02903_ _02908_ _02745_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08056__A1 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10337__B _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06067__B1 _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ _01181_ _01324_ _01454_ _02001_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_15_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08093_ as2650.indirect_target\[9\] _02757_ _02842_ _02844_ _02845_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_43_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07044_ net193 _01773_ _01782_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08995_ _03686_ _03650_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ _01319_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06790__A1 _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input27_I bus_in_timers[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07877_ _01721_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_108_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_3_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__B _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09616_ _02943_ _04301_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06828_ _01204_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06776__I _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06759_ _01674_ _01627_ _01680_ net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_09547_ _04232_ _03634_ _02468_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_1422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_65_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09478_ _04084_ _04086_ _04163_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_136_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08429_ _00649_ _03123_ _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11440_ _00224_ clknet_leaf_37_wb_clk_i as2650.ivectors_base\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11371_ _00167_ clknet_leaf_70_wb_clk_i net233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ _04825_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11857__I net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10253_ _04830_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_123_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10184_ _04697_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09562__A4 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08770__A2 _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_135_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_135_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06686__I _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06619__C _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10001__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11707_ _00491_ clknet_leaf_22_wb_clk_i as2650.stack\[6\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11638_ _00422_ clknet_leaf_13_wb_clk_i as2650.stack\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09786__A1 _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11569_ _00353_ clknet_leaf_41_wb_clk_i as2650.stack\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09538__A1 _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08210__A1 _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _02559_ _02562_ _02568_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09681__B _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08780_ _01506_ _03457_ _03458_ _03476_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05992_ net222 _00976_ _00992_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07731_ _02499_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07662_ net392 _02340_ _02434_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06524__A1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10320__A2 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09401_ _04084_ _04086_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06613_ as2650.debug_psl\[0\] _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07593_ _02373_ _02383_ _02386_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_1618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _01499_ _01017_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06544_ _00827_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09263_ _01022_ _00887_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06475_ _01437_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08214_ _02951_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08029__A1 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09194_ _00716_ _00873_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08145_ as2650.instruction_args_latch\[13\] _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_112_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08076_ _02800_ _01845_ _02817_ _02816_ _02828_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_82_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06460__B1 _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07027_ _01934_ _01935_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_25_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05675__I as2650.debug_psl\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08201__A1 _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07004__A2 _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08201__B2 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold23 _02308_ net367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08978_ _03617_ _03618_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xhold34 _02369_ net378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__06763__A1 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold45 net445 net389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07960__B1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold56 net95 net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold67 _02068_ net411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07929_ _01251_ _01333_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold78 net451 net422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output133_I net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold89 wbs_dat_i[4] net435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08504__A2 _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10940_ _05375_ _05297_ _05298_ _00763_ _05376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06515__A1 _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06515__B2 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10311__A2 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ _05262_ _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_119_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08654__C _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09768__A1 _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _00207_ clknet_leaf_68_wb_clk_i as2650.instruction_args_latch\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11354_ _00150_ clknet_leaf_108_wb_clk_i wb_counter\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10305_ _04224_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10491__I _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11285_ _00081_ clknet_leaf_142_wb_clk_i net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_56_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10236_ _01238_ _02917_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_52_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09940__A1 net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08743__A2 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _04705_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06754__A1 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08829__C _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10098_ as2650.stack\[3\]\[9\] _04682_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07305__I _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06809__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_32_wb_clk_i clknet_4_6__leaf_wb_clk_i clknet_leaf_32_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_152_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06260_ _01232_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_26_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06191_ _01148_ _01149_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07234__A2 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09950_ _01477_ _04428_ _04585_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__05796__A2 _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06993__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ _01419_ _01212_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_146_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09881_ as2650.stack\[5\]\[9\] _04540_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_146_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A2 _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08832_ _03523_ _03524_ _03525_ _03526_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06745__A1 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10541__A2 _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05975_ _00943_ _00977_ _00956_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08763_ _01879_ _03459_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_139_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07714_ _02482_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08498__A1 as2650.stack\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08694_ _03374_ _03391_ _03393_ _03344_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08498__B2 as2650.stack\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_101_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07645_ wb_counter\[25\] _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_62_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07576_ _02358_ _02371_ _02372_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_152_1497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05720__A2 _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06527_ _01241_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09315_ _03997_ _03999_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06458_ _01344_ _01361_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09246_ _00826_ _03931_ _01498_ _00913_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_88_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09177_ _01569_ _02576_ _02591_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_135_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06389_ _00844_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ _02788_ _01920_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ _02812_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_92_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06984__A1 _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output250_I net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11070_ _04769_ _05142_ _04721_ _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_124_1599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput102 net393 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10021_ _04629_ _04625_ _04630_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06736__A1 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10923_ _05295_ _05350_ _05360_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06964__I as2650.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10854_ _05294_ _05295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_1672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10785_ as2650.stack\[6\]\[4\] _05238_ _05239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_136_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07795__I _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11406_ _00190_ clknet_leaf_45_wb_clk_i as2650.indirect_target\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08964__A2 _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11337_ _00133_ clknet_leaf_145_wb_clk_i wb_counter\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_150_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_150_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_162_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11268_ _00064_ clknet_leaf_137_wb_clk_i net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_10219_ _01372_ _04796_ _04737_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_11199_ as2650.stack\[9\]\[7\] _05557_ _05561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_145_Left_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05760_ _00688_ _00752_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09677__B1 _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05950__A2 _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07035__I _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05691_ _00704_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09692__A3 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07430_ _01943_ _02147_ _02148_ _02258_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_114_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06874__I _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_122_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07361_ _02118_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06312_ _01282_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_84_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09100_ _03722_ _03789_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07292_ _02130_ _02135_ _02138_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08652__B2 as2650.stack\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_154_Left_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09031_ _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06243_ _01215_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_147_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06174_ _01079_ _01145_ _01146_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__08404__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05769__A2 _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09933_ net142 _01466_ _04572_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06114__I _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09864_ _01777_ _04526_ _04531_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_163_Left_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08815_ _03190_ _01909_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_77_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09795_ _01681_ _03142_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_20_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08746_ _01865_ _03375_ _03443_ _03197_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_169_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05958_ _00744_ as2650.instruction_args_latch\[12\] _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10278__A1 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08677_ as2650.stack\[0\]\[5\] _02491_ _02498_ as2650.stack\[1\]\[5\] _03130_ _03377_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_85_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05889_ _00800_ as2650.regs\[4\]\[2\] _00894_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_85_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _02407_ _02413_ _02414_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07694__A2 _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07559_ wb_counter\[8\] _02354_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_81_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10570_ _05098_ _05095_ _05099_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_146_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ _03914_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10202__A1 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11122_ _05465_ _05508_ _05512_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06024__I _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11053_ as2650.stack\[0\]\[11\] _05461_ _05468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06709__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10004_ as2650.stack\[4\]\[13\] _04616_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09659__B1 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09123__A2 _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10906_ _05320_ _05343_ _05344_ _05345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08882__A1 _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10837_ _04440_ _02559_ _05279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_66_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11105__I _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08634__A1 _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ as2650.regs\[6\]\[7\] _05227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10441__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05999__A2 as2650.cycle\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10699_ _05174_ _05184_ _05185_ _00908_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_144_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09954__B _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10744__A2 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_143_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06930_ _01844_ _01827_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_input1_I bus_in_gpios[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__A2 _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06861_ as2650.debug_psl\[3\] _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08600_ _02497_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05812_ as2650.regs\[0\]\[3\] _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06792_ _01712_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09580_ _01855_ _03744_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09114__A2 _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08531_ _03102_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05743_ _00754_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05674_ _00663_ _00686_ _00687_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08462_ _01546_ _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06479__A3 _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07413_ _02115_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08393_ as2650.stack\[11\]\[14\] _02510_ _02513_ as2650.stack\[10\]\[14\] _03114_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11015__I _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07344_ _02183_ _01772_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07428__A2 _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07275_ net131 _02119_ _02122_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06226_ _01195_ _01198_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09014_ _03580_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06157_ _01129_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_108_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold120 wbs_stb_i net466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_143_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09050__A1 _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input57_I ram_bus_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06088_ _01065_ _01066_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_74_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _04563_ net151 _04564_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10499__A1 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _04519_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_126_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_126_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07364__A1 _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08561__B1 _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09778_ _04431_ _04457_ _04460_ _01454_ _04445_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_119_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09105__A2 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08729_ _01865_ _03280_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output213_I net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _00524_ clknet_leaf_133_wb_clk_i as2650.stack\[0\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08864__A1 _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11671_ _00455_ clknet_leaf_98_wb_clk_i as2650.regs\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10622_ as2650.stack\[7\]\[11\] _05130_ _05134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06019__I _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10423__A1 _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10553_ _05084_ _05085_ _05087_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06463__B _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10974__A2 _05286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08234__I _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _04659_ _05038_ _05041_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05602__B2 as2650.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11105_ _05494_ _05502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_104_1767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11036_ as2650.stack\[0\]\[6\] _05451_ _05456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07355__A1 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08855__A1 _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08607__A1 _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10414__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08083__A2 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__I1 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07060_ _01964_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_11_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06011_ _01009_ net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_140_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput203 net203 la_data_out[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05841__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput214 net214 la_data_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput225 net225 last_addr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_65_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput236 net236 last_addr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07983__I _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput247 net247 requested_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_122_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput258 net258 rom_bus_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput269 net269 wbs_dat_o[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06397__A2 _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_166_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08791__B1 _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07962_ as2650.irqs_latch\[2\] as2650.irqs_latch\[3\] _02720_ _02721_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09701_ net1 net9 net25 net17 _04383_ _04384_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_103_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06913_ _01827_ _01828_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07893_ _01332_ _01304_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_120_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08543__B1 _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09632_ _01754_ _01886_ _02578_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06844_ _01719_ _01762_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_121_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10849__I _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09099__A1 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09563_ _03847_ _04248_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_155_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06775_ _01695_ _01100_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_72_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08514_ _02554_ _02555_ _03218_ _01219_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_05726_ _00601_ net430 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_91_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09494_ _04164_ _04166_ _04167_ _04179_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__07223__I _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07113__A4 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08445_ _02665_ _02943_ _03161_ _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_05657_ _00670_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_108_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05588_ as2650.PC\[3\] _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08376_ _03020_ _03097_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_129_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07327_ net137 _02168_ _02150_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05678__I _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06085__A1 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08054__I _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07258_ _01553_ _02083_ _02105_ _02106_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_1734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_76_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06209_ _01130_ _01172_ _01181_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07189_ net91 net108 _02046_ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_128_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08657__C _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06560__A2 _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08837__A1 _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11723_ _00507_ clknet_leaf_76_wb_clk_i as2650.regs\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11654_ _00438_ clknet_leaf_93_wb_clk_i as2650.regs\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10605_ _05117_ _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11585_ _00369_ clknet_leaf_93_wb_clk_i as2650.regs\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05588__I as2650.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ _05072_ _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_150_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10467_ as2650.stack\[2\]\[7\] _05027_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10398_ _01557_ _01383_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08773__B1 _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11019_ as2650.stack\[0\]\[1\] _05441_ _05444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07879__A2 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10883__A1 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10669__I _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06560_ _01154_ _01505_ _01514_ net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__07043__I net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10635__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06491_ _01453_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07500__A1 net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07978__I _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08230_ _02904_ _02964_ _02965_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08161_ as2650.indirect_target\[14\] _02904_ _02713_ _02907_ _02718_ _02908_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_28_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07112_ _02000_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06067__B2 _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08092_ _01258_ _02843_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_126_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07043_ net306 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05814__A1 _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08994_ _03598_ _03599_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07945_ _02616_ _02644_ _02703_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07876_ _01326_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_108_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09615_ _04294_ _04295_ _04298_ _04299_ _04300_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_39_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10579__I _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06827_ _00872_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09546_ _03635_ _03662_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06758_ net253 _01527_ _01531_ _01679_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_65_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05709_ _00721_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_09477_ _03981_ _04082_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06689_ _01078_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06792__I _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08428_ _03107_ _03065_ _03146_ _03061_ _03147_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_163_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08359_ _02614_ _03075_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_151_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11370_ _00166_ clknet_leaf_70_wb_clk_i net232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_145_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09795__A2 _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _04360_ _04818_ _04896_ _04814_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_131_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10252_ _01084_ _04696_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05820__A4 _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10183_ _02659_ _04728_ _04759_ _04760_ _04761_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_121_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10865__A1 _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_104_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_104_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11706_ _00490_ clknet_leaf_40_wb_clk_i as2650.stack\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08038__A2 _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11637_ _00421_ clknet_leaf_11_wb_clk_i as2650.stack\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11568_ _00352_ clknet_leaf_41_wb_clk_i as2650.stack\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08850__C _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10519_ _04651_ _05059_ _05063_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11499_ _00283_ clknet_leaf_125_wb_clk_i as2650.stack\[5\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08422__I _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06221__A1 _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05991_ _00982_ _00983_ _00975_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_100_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07730_ _02498_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07661_ wb_counter\[29\] _02440_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_117_1722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06524__A2 _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09400_ _03973_ _03979_ _04085_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06612_ wb_debug_carry _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_137_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ net402 _02376_ _02385_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_103_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09331_ _04012_ _04016_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_157_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06543_ _01500_ net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_146_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06288__A1 _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09262_ _03946_ _03947_ _03875_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_145_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06474_ _01436_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08213_ _01332_ _01308_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09193_ _00754_ _00896_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08144_ _02632_ _02891_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08075_ _02827_ _01864_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_rebuffer12_I _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06460__A1 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07026_ _01915_ _01918_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09529__A2 _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08737__B1 _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold13 net435 net357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08977_ _03625_ _03666_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_122_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold24 _00123_ net368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_157_1513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold35 _00140_ net379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08488__B _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold46 net100 net390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_2_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07928_ as2650.indirect_target\[1\] _02680_ _02687_ _01453_ _02688_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xhold57 net452 net401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold68 net447 net412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold79 net465 net423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07859_ _01534_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output126_I net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07712__A1 _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10870_ _04247_ _05302_ _05310_ _05311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09529_ _03684_ _03773_ _03776_ _03600_ _04214_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_116_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09217__A1 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11422_ _00206_ clknet_leaf_64_wb_clk_i as2650.instruction_args_latch\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06027__I _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10772__I _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11353_ _00149_ clknet_leaf_108_wb_clk_i wb_counter\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05866__I _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ as2650.regs\[5\]\[3\] _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_120_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11284_ _00080_ clknet_leaf_139_wb_clk_i net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_56_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_56_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10235_ _04247_ _04729_ _04792_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_52_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold28_I wbs_dat_i[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10166_ _04731_ _04741_ _04743_ _04744_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_7_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06754__A2 _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10097_ _04645_ _04681_ _04683_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_112_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08845__C _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10999_ _05369_ _05398_ _05426_ _05427_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_31_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10066__A2 _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08417__I _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06809__A3 _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06690__A1 net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06190_ _01162_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_160_Right_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_72_wb_clk_i clknet_4_15__leaf_wb_clk_i clknet_leaf_72_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_108_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08900_ _03582_ _03591_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_111_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09880_ _01883_ _04539_ _04541_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_146_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07991__I _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ as2650.stack\[15\]\[10\] _03466_ _03246_ as2650.stack\[14\]\[10\] _03520_
+ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__06745__A2 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07942__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_151_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08762_ _00592_ _03441_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05974_ _00973_ _00939_ _00975_ _00976_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_105_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07713_ _01274_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_159_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08693_ _02776_ _03108_ _03228_ _03392_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08498__A2 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11018__I _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07644_ _02423_ _02425_ _02427_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_152_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07575_ net388 _02361_ _02368_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05720__A3 _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ _03997_ _03999_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_1584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06526_ _01477_ as2650.cycle\[8\] _01486_ _01247_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_146_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09245_ _00816_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06457_ _01419_ _01378_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_88_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11006__A1 _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09176_ _01570_ _03714_ _03860_ _03862_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_135_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06388_ _01350_ _01351_ _01352_ _00872_ _00736_ _00706_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_135_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _02866_ _02876_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06433__A1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08058_ net65 _02763_ _02811_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_109_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07009_ _01915_ _01918_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10020_ as2650.stack\[10\]\[1\] _04627_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output243_I net243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09922__A2 net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput103 net403 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06736__A2 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06310__I _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09686__A1 as2650.cycle\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10922_ as2650.regs\[4\]\[4\] _05335_ _05359_ _05294_ _05360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10853_ _03816_ _05259_ _05294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_116_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10784_ _05231_ _05238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f__01549_ clknet_0__01549_ clknet_1_0__leaf__01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11405_ _00189_ clknet_leaf_45_wb_clk_i as2650.indirect_target\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09610__A1 _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11336_ _00132_ clknet_leaf_145_wb_clk_i wb_counter\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11267_ _00063_ clknet_leaf_135_wb_clk_i net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_10218_ _01503_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11198_ _05455_ _05556_ _05560_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06727__A2 _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10149_ _04727_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_141_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10170__C _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07316__I _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05950__A3 _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05690_ _00703_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_153_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10677__I _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__I _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ _02191_ _02196_ _02198_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06311_ _01281_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10444__C1 _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ net292 _02137_ _02128_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_1555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07986__I _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09030_ _03721_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06890__I _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06242_ _01214_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold117_I wbs_dat_i[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06173_ net64 _01079_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09601__A1 _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_130_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09932_ _02677_ _04570_ _04574_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07215__I0 net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ as2650.stack\[5\]\[2\] _04528_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06718__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08814_ _03343_ _01909_ _03192_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09794_ _01526_ _04474_ _04475_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08745_ _03312_ _03440_ _03442_ _01445_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05957_ _00630_ _00632_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09668__A1 _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07670__B _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08676_ as2650.stack\[3\]\[5\] _01691_ _01967_ as2650.stack\[2\]\[5\] _03376_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05888_ _00689_ _00893_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_132_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A1 _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ net86 _02410_ _02401_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07558_ _02357_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_81_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06509_ _01089_ _01316_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09840__A1 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07489_ _01553_ _02059_ _02304_ _02063_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_8_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07896__I _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09228_ _00728_ _00775_ _01012_ _01014_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_49_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output193_I net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ _03838_ _03840_ _03845_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_121_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11211__I _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06305__I _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11121_ as2650.stack\[14\]\[10\] _05509_ _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08159__A1 _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11052_ _01927_ _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06709__A2 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10003_ _01940_ _04615_ _04617_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_34_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07136__I _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06040__I _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09659__B2 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06975__I _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10905_ _04310_ _05312_ _05344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold95_I wbs_dat_i[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06893__A1 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ _03706_ _02580_ _05278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10767_ _05178_ _05222_ _05223_ _05226_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_82_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09831__A1 as2650.debug_psu\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07842__B1 _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10698_ _05182_ _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11319_ _00115_ clknet_leaf_104_wb_clk_i net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_129_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06860_ _01716_ _01777_ _01778_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05811_ _00820_ net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06791_ _01697_ _01701_ _01711_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08530_ _03103_ _03189_ _03233_ _03234_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_145_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05742_ as2650.regs\[1\]\[6\] as2650.regs\[5\]\[6\] _00753_ _00754_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08322__B2 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _01355_ _03171_ _03173_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05673_ as2650.insin\[0\] _00663_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08873__A2 _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07412_ _02237_ _02243_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11209__A1 as2650.stack\[9\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ _03109_ _03110_ _03111_ _03112_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10417__C1 _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07343_ _02141_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08625__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10432__A2 _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_147_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _03704_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06225_ _01197_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_131_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold110 wbs_dat_i[30] net456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06156_ _01103_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold121 wbs_dat_i[22] net467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06087_ _00810_ _00931_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_74_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05611__A2 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09915_ _03174_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09846_ net47 as2650.irqs_latch\[5\] _04514_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_126_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07364__A2 _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_87_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _04439_ _03761_ _04458_ _04459_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_06989_ _01871_ _01899_ _01900_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08728_ _03398_ _03423_ _03426_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06795__I _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08313__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09171__I _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output206_I net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ as2650.stack\[15\]\[4\] _01691_ _01967_ as2650.stack\[14\]\[4\] _02519_ _03360_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_1_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A1 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11670_ _00454_ clknet_leaf_98_wb_clk_i as2650.regs\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10621_ _05100_ _05129_ _05133_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_27_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09813__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_22_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10552_ as2650.stack\[15\]\[4\] _05086_ _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ as2650.stack\[2\]\[13\] _05039_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_129_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_129_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06035__I _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07052__A1 as2650.page_reg\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__B _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05874__I _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11104_ _05447_ _05495_ _05501_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11035_ _01852_ _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07107__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11116__I _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06866__A1 _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10819_ _05260_ _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11799_ _00578_ clknet_leaf_28_wb_clk_i as2650.stack\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09804__B2 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06618__A1 as2650.insin\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06094__A2 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07291__A1 net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06010_ _00956_ _00964_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09568__B1 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput204 net204 la_data_out[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput215 net215 la_data_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_3_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09032__A2 _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput226 net226 last_addr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput237 net237 le_hi_act vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_65_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10690__I _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput248 net248 requested_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput259 net259 rom_bus_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07961_ as2650.irqs_latch\[4\] as2650.irqs_latch\[5\] _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_26_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09700_ net5 net13 net29 net21 _01518_ _01520_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_06912_ _01812_ _01814_ _01826_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07892_ _02653_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09631_ _02813_ _04313_ _04316_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06843_ as2650.PC\[1\] _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10350__A1 _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09562_ _04224_ _04231_ _04239_ _04247_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_121_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06774_ _01236_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_151_1508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08513_ _03213_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_52_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05725_ _00714_ _00737_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_91_1654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09493_ _04168_ _04169_ _04178_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_66_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06857__A1 _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08444_ _03158_ _03159_ _02579_ _03160_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_93_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05656_ net227 net226 _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_59_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08375_ as2650.instruction_args_latch\[9\] as2650.instruction_args_latch\[10\] _03096_
+ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_163_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05587_ _00592_ _00597_ _00600_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_119_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07326_ _02117_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_22_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06085__A2 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07257_ _02086_ net130 _02087_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09559__B1 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06208_ _01180_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_76_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07188_ _02049_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06139_ net60 _01111_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_112_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output156_I net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10105__I _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08534__A1 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09829_ _01857_ _02485_ _04506_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07842__C _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10341__A1 _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06560__A3 _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11722_ _00506_ clknet_leaf_77_wb_clk_i as2650.regs\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06848__A1 _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11653_ _00437_ clknet_leaf_92_wb_clk_i as2650.regs\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10604_ _05115_ _05123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11584_ _00368_ clknet_leaf_93_wb_clk_i as2650.regs\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10535_ _05073_ _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_145_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold58_I net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10466_ _04641_ _05026_ _05030_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10397_ _04733_ _04968_ _04969_ _04740_ _01837_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_23_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05587__A1 _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_97_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_97_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_161_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11018_ _01759_ _05443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_wb_clk_i clknet_4_6__leaf_wb_clk_i clknet_leaf_26_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08828__A2 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__B _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06839__A1 _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06490_ _01452_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07500__A2 _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10685__I _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_4_13__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08160_ _02905_ _01298_ _02678_ _02906_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_32_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07111_ _01472_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08091_ _02644_ _02634_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_144_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07042_ as2650.page_reg\[1\] _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_168_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09005__A2 _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07016__A1 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06403__I _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08993_ _03680_ _03681_ _03684_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07944_ _02702_ _02701_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08516__A1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07875_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10323__A1 _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06559__B _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09614_ _01576_ _02470_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06826_ _00606_ _01741_ _01745_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_69_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_69_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09545_ _03670_ _03842_ _04226_ _04230_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_151_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06757_ _01675_ _01678_ _01078_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_78_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05708_ _00720_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09476_ _04125_ _04161_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10626__A2 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06688_ _01615_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_66_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08427_ _00644_ _03061_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05639_ as2650.page_reg\[1\] _00646_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10595__I _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05689__I _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08358_ _02601_ _00844_ _01437_ _03079_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_78_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09244__A2 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07309_ net294 _02137_ _02128_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08289_ _02761_ _03015_ _03016_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _01399_ _04820_ _04895_ _04819_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_81_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07837__C _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10251_ _04382_ _04761_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_30_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08755__A1 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10182_ _04707_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10562__A1 _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07853__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08507__A1 _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11705_ _00489_ clknet_leaf_40_wb_clk_i as2650.stack\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11465__CLK clknet_4_12__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_144_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_144_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11636_ _00420_ clknet_leaf_11_wb_clk_i as2650.stack\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_1442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06049__A2 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11567_ _00351_ clknet_leaf_12_wb_clk_i as2650.stack\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08994__A1 _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07797__A2 _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10518_ as2650.stack\[1\]\[10\] _05060_ _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11498_ _00282_ clknet_leaf_137_wb_clk_i as2650.stack\[5\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10449_ _05017_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_163_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07319__I _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08746__A1 _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10553__A1 _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06221__A2 _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05990_ _00980_ net255 _00989_ _00990_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA_clkbuf_leaf_141_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07660_ _02439_ _02436_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06611_ net304 _01554_ _01555_ net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_149_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07591_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_103_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09330_ _04013_ _04014_ _04015_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_157_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06542_ _01499_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_157_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06288__A2 _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07485__A1 _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09261_ _00716_ _00854_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06473_ _01192_ _01197_ _01189_ _01217_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_111_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08212_ _01485_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09192_ _03875_ _03876_ _03877_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08143_ _02889_ _02890_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07237__A1 _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08074_ _02786_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_31_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05799__A1 _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__A1 _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07025_ as2650.PC\[12\] _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_105_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07229__I _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08737__B2 as2650.stack\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold14 net98 net358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_08976_ _03664_ _03665_ _03667_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input32_I bus_in_timers[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold25 net431 net369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold36 net462 net380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07960__A2 _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold47 net438 net391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07927_ _02000_ _02686_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xhold58 net78 net402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold69 net449 net413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09162__A1 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07858_ _02611_ _02621_ _02622_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06809_ _01727_ _01509_ _01699_ _01729_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_39_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output119_I net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07789_ net216 _02485_ _02478_ _02553_ _02557_ _01462_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_0_151_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07899__I _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09528_ _01283_ _03682_ _03603_ _02920_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_78_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07476__A1 net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _04140_ _04141_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09217__A2 net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11421_ _00205_ clknet_leaf_62_wb_clk_i as2650.instruction_args_latch\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11352_ _00148_ clknet_leaf_108_wb_clk_i wb_counter\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10303_ _04841_ _04789_ _04874_ _04835_ _04879_ _04840_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__06451__A2 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11283_ _00079_ clknet_leaf_107_wb_clk_i net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_56_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10234_ _01599_ _04793_ _04807_ _04809_ _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_123_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_5_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06203__A2 _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _04718_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06978__I as2650.PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05882__I _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05962__A1 _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10096_ as2650.stack\[3\]\[8\] _04682_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09153__A1 _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07703__A2 _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08900__A1 _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10998_ as2650.regs\[0\]\[5\] _05405_ _05427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07602__I _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09700__I0 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10963__I _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11619_ _00403_ clknet_leaf_18_wb_clk_i as2650.stack\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08967__A1 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08719__A1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_41_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_41_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_123_1771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ as2650.stack\[12\]\[10\] _02526_ _02529_ as2650.stack\[13\]\[10\] _03525_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06888__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07942__A2 _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08761_ _02825_ _03288_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05973_ _00954_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_105_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07712_ _01943_ _02480_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_159_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08692_ _03229_ _01830_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07643_ net89 _02426_ _02418_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_101_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_101_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_4_3__f_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07574_ wb_counter\[12\] _02370_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_117_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07512__I _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09447__A2 _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09313_ _03942_ _03998_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06525_ _01479_ _01484_ _01485_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07458__A1 net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09244_ _01027_ _00888_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06456_ _00769_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06128__I _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08771__C _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09175_ _01336_ _01222_ _01337_ _03861_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__11006__A2 _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06387_ net196 _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_135_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08126_ as2650.ivectors_base\[7\] _02852_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_96_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08057_ _01153_ _01136_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_92_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07008_ _01917_ _01906_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08186__A2 _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput104 net466 net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output236_I net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ _03600_ _03650_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08011__C _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09135__A1 _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09686__A2 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10921_ _04324_ _05263_ _05358_ _05359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_54_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10852_ _05261_ _05282_ _05289_ _05293_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_135_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10783_ _05229_ _05237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_45_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06038__I _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10783__I _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08949__A1 _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _00188_ clknet_leaf_46_wb_clk_i as2650.indirect_target\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_105_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__A2 as2650.debug_psl\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_1722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11335_ _00131_ clknet_leaf_153_wb_clk_i wb_counter\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11266_ _00062_ clknet_leaf_134_wb_clk_i net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__10508__A1 as2650.stack\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10217_ _04732_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11653__CLK clknet_leaf_92_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11197_ as2650.stack\[9\]\[6\] _05557_ _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10148_ _04706_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_141_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09126__A1 _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10079_ _04629_ _04668_ _04672_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07688__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05950__A4 _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_59_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06360__A1 _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06310_ _01280_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10444__B1 _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07290_ _02136_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06241_ _01213_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06172_ net35 _01133_ _01144_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_131_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09601__A2 _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07612__A1 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_68_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_145_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09931_ net141 _01466_ _04572_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07215__I1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _01760_ _04526_ _04530_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07507__I as2650.wb_hidden_rom_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08813_ _02861_ _03507_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09793_ _02573_ _01706_ _04465_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__11029__I _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05956_ _00957_ _00959_ _00960_ _00590_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_139_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08744_ _00592_ _03441_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09668__A2 _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_77_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_1674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07679__A1 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ _03243_ _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_124_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08876__B1 _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05887_ as2650.regs\[0\]\[2\] _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07626_ wb_counter\[22\] _02412_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_85_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07557_ _02319_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_81_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_137_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06508_ _01468_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_107_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ net94 _02058_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_98_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06439_ _01401_ _01359_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_40_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09227_ _00775_ _01012_ _01014_ _00729_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09158_ _03679_ _03841_ _03842_ _03844_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_72_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output186_I net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08109_ as2650.indirect_target\[10\] _02680_ _02844_ _02859_ _02860_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_20_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08800__B1 _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09089_ _01169_ _03771_ _03773_ _03694_ _03778_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_114_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11120_ _05463_ _05508_ _05511_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08159__A2 _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11051_ _05465_ _05460_ _05466_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11163__A1 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10002_ as2650.stack\[4\]\[12\] _04616_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_95_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09659__A2 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10904_ _04224_ _05302_ _05342_ _05343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11218__A2 _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10835_ _05274_ _04725_ _05276_ _05277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08095__A1 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold88_I wbs_dat_i[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10766_ as2650.regs\[6\]\[6\] _05226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10977__A1 _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09831__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__B2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ _05180_ _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_129_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09079__I _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11318_ _00114_ clknet_leaf_105_wb_clk_i net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_143_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11249_ _00045_ clknet_leaf_125_wb_clk_i as2650.stack\[11\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09898__A2 _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05810_ _00796_ _00818_ _00819_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06790_ _01505_ _01707_ _01708_ _01710_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__06581__A1 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05741_ as2650.debug_psl\[4\] _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_136_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08322__A2 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08460_ as2650.ivectors_base\[4\] _03172_ _03167_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05672_ _00681_ _00685_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08158__I _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07062__I _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07411_ net276 _02238_ _02242_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08391_ as2650.stack\[4\]\[14\] _02493_ _02500_ as2650.stack\[5\]\[14\] _02521_ _03112_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_114_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07342_ net124 _02139_ _02175_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10417__B1 _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08086__A1 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07833__A1 _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ _02120_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09012_ _02466_ _02587_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06224_ _01196_ _01151_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_104_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06406__I net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold100 wbs_dat_i[21] net446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09586__A1 _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06155_ _01116_ _01127_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold111 wbs_dat_i[5] net457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__09050__A3 _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06086_ net349 _00930_ _00933_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_1505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09914_ as2650.cycle\[1\] _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05611__A3 _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08010__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09845_ _04518_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_126_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08561__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07681__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _01268_ _04450_ _04429_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06988_ as2650.stack\[12\]\[9\] _01884_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08727_ _02670_ _03425_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05939_ _00748_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_69_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09510__A1 _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08658_ as2650.stack\[12\]\[4\] _03305_ _03306_ as2650.stack\[13\]\[4\] _03359_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_96_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10120__A2 _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ wb_counter\[17\] wb_counter\[18\] _02392_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_83_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08589_ _02490_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10620_ as2650.stack\[7\]\[10\] _05130_ _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10551_ _05075_ _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07824__A1 _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10482_ _04655_ _05038_ _05040_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09577__A1 _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08531__I _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07052__A2 _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11103_ as2650.stack\[14\]\[3\] _05497_ _05501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09329__A1 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11034_ _05453_ _05450_ _05454_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06051__I _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05890__I _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09501__A1 _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__A1 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10111__A2 _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08068__A1 _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10818_ _03817_ _05259_ _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11798_ _00577_ clknet_leaf_25_wb_clk_i as2650.stack\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06618__A2 _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10749_ _05214_ _05215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__A1 _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09568__B2 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10178__A2 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput205 net205 la_data_out[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput216 net216 la_data_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput227 net227 last_addr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput238 net238 le_lo_act vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput249 net249 requested_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_166_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07960_ as2650.indirect_target\[2\] _01259_ _02713_ _02717_ _02718_ _02719_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06911_ as2650.PC\[4\] _01826_ _01814_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07891_ _01294_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_120_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_155_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09740__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08543__A2 _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ _02615_ _04314_ _04315_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06842_ _01716_ _01760_ _01761_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06554__A1 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09561_ _01168_ _04240_ _04246_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_121_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_97_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06773_ _01693_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05724_ _00706_ _00722_ _00731_ _00736_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_91_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08512_ _02639_ _03216_ _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09492_ _04171_ _04173_ _04174_ _04177_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_72_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05655_ _00668_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08443_ _01216_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_72_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _03068_ _03095_ _02999_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05586_ as2650.indirect_target\[7\] _00599_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07325_ _02162_ _02165_ _02167_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07806__A1 net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11042__I _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07256_ _02084_ net161 _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06207_ _01173_ _01179_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_76_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07187_ net90 net107 _02046_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10169__A2 _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input62_I rom_bus_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06138_ _00665_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06069_ net221 _01050_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11118__A1 _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output149_I net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09828_ _04449_ _03754_ _03146_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_154_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09759_ _01704_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _00505_ clknet_leaf_82_wb_clk_i as2650.regs\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11652_ _00436_ clknet_leaf_92_wb_clk_i as2650.regs\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10603_ _05082_ _05116_ _05122_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_61_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09798__A1 _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11583_ _00367_ clknet_leaf_91_wb_clk_i as2650.regs\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10534_ _05072_ _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07586__B _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10465_ as2650.stack\[2\]\[6\] _05027_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08261__I _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10396_ _03856_ _01504_ _04734_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_62_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08773__A2 _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05587__A2 _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10580__A2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_131_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08525__A2 _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11017_ _05436_ _05439_ _05442_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_1775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08289__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_66_wb_clk_i clknet_4_13__leaf_wb_clk_i clknet_leaf_66_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09789__A1 _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07110_ _01998_ _01266_ _01469_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_126_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08090_ _02838_ _02841_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_67_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08461__A1 _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09695__C _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07041_ _01930_ _01947_ _01948_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_168_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05795__I _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08213__A1 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09961__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08992_ _03683_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_23_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07943_ _02642_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08516__A2 _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07874_ _01506_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_3_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09613_ _01564_ _03720_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_108_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06825_ _01742_ _01744_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09544_ _03672_ _03841_ _04227_ _02468_ _04229_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_06756_ _01543_ _01677_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08774__C _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05707_ _00719_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09475_ _03928_ _04089_ _04127_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06687_ _01614_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08426_ _03135_ _03145_ _02552_ _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05638_ as2650.instruction_args_latch\[14\] _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_110_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ _02675_ _03078_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_78_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07308_ _02114_ wb_counter\[6\] _02152_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08452__A1 as2650.ivectors_base\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08288_ _03006_ _01315_ _02861_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_127_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07239_ _02066_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10250_ _02677_ _04728_ _04761_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08204__A1 _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output266_I net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10181_ _01412_ _04712_ _04727_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10562__A2 _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08684__C _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11704_ _00488_ clknet_leaf_13_wb_clk_i as2650.stack\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11635_ _00419_ clknet_leaf_10_wb_clk_i as2650.stack\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11566_ _00350_ clknet_leaf_13_wb_clk_i as2650.stack\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10250__A1 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _04649_ _05059_ _05062_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11497_ _00281_ clknet_leaf_127_wb_clk_i as2650.stack\[5\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_1508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10448_ _05018_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_150_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_163_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09943__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10379_ _01385_ _04820_ _04952_ _04817_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_81_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10553__A2 _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06509__A1 _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06610_ web_behavior\[1\] _01553_ clknet_leaf_149_wb_clk_i _01555_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07590_ _02073_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06541_ _01498_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06472_ _01192_ _01434_ _01189_ _01322_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09260_ _00754_ _00873_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07070__I _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ _02623_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09191_ _00717_ _00755_ _00874_ _00855_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_28_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08142_ _02636_ _00958_ _01708_ _02794_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07237__A2 net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08073_ _01147_ _02825_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05799__A2 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06996__A1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07024_ _00915_ _01753_ _01932_ _01734_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_144_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09934__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08737__A2 _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10544__A2 _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _03637_ _03666_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold15 _02311_ net359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_122_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold26 _02316_ net370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold37 net80 net381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07926_ _01326_ _02682_ _02685_ _01319_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xhold48 net93 net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_157_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold59 net442 net403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_1661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input25_I bus_in_timers[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09162__A2 _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07857_ _02003_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06808_ _01728_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07788_ _02556_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09527_ _03823_ _04200_ _04212_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_151_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06739_ net251 _01617_ _01531_ _01662_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_116_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07476__A2 _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09458_ _04128_ _04131_ _04143_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_149_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08409_ as2650.stack\[3\]\[15\] _02510_ _02513_ as2650.stack\[2\]\[15\] _03129_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_137_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09389_ _04061_ _04063_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_93_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11420_ _00204_ clknet_leaf_64_wb_clk_i as2650.instruction_args_latch\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_43_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10232__A1 _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _00147_ clknet_leaf_108_wb_clk_i wb_counter\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10302_ _04877_ _04878_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06324__I _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11282_ _00078_ clknet_leaf_107_wb_clk_i net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_132_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09925__A1 _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10233_ _04810_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06739__A1 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08679__C _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _01615_ _04742_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_140_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10095_ _04669_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06994__I as2650.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06911__A1 as2650.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10997_ _05424_ _05425_ _05397_ _05426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09700__I1 net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08664__A1 _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_106_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_152_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11618_ _00402_ clknet_leaf_23_wb_clk_i as2650.stack\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11549_ _00333_ clknet_leaf_8_wb_clk_i as2650.stack\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10526__A2 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_115_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08760_ _03226_ _03455_ _03456_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05972_ _00947_ _00974_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_139_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07065__I _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_81_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_81_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_105_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07711_ _02464_ _02479_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08691_ _01831_ _03283_ _03390_ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_10_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07642_ _02339_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_101_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07573_ wb_counter\[11\] _02364_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11462__D _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09312_ _03939_ _03943_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06524_ _01480_ _01305_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06409__I _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08655__A1 _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09243_ _00728_ _01020_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06455_ _01344_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_1649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06386_ _00865_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09174_ net216 _03722_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06418__B1 _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08125_ _02837_ _02872_ _02873_ _02874_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_47_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06969__A1 _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08056_ _02611_ _02808_ _02810_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_109_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07007_ _01905_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_101_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput105 net428 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_122_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11190__A2 _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08958_ _03602_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05944__A2 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09135__A2 _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output131_I net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _02669_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08889_ _01343_ _01227_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10920_ _05320_ _05357_ _05358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10851_ _05292_ _05260_ _05293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10782_ _05082_ _05230_ _05236_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_45_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10205__A1 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11403_ _00187_ clknet_leaf_44_wb_clk_i as2650.indirect_target\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09610__A3 _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11334_ _00130_ clknet_leaf_154_wb_clk_i wb_counter\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05632__A1 _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _00061_ clknet_leaf_134_wb_clk_i net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_103_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold33_I net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10216_ _01194_ _02469_ _01696_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_120_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _05453_ _05556_ _05559_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_145_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10147_ _04697_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_141_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10078_ as2650.stack\[3\]\[1\] _04670_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07688__A2 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06240_ _01212_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_1557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06171_ _01143_ _01132_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_130_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05623__A1 _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09930_ _02659_ _04570_ _04573_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06899__I _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09861_ as2650.stack\[5\]\[1\] _04528_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08812_ _02846_ _03096_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10214__I _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09792_ _04431_ _04470_ _04473_ _01454_ _04445_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05926__A2 _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08743_ _01826_ _01848_ _03387_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05955_ _00633_ _00637_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09668__A3 _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07679__A2 net238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _03224_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_1795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05886_ _00892_ net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_132_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07625_ wb_counter\[20\] wb_counter\[21\] _02404_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_85_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07556_ _02341_ _02355_ _02356_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10435__A1 _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_137_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06507_ _01264_ _01304_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_137_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07487_ _02097_ _02059_ _02303_ _02063_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_14_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_98_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05978__I net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09226_ _03890_ _03900_ _03911_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06438_ _00828_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09157_ _03646_ _03647_ _03843_ _01231_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_115_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06369_ _01332_ _01333_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_EDGE_ROW_141_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08108_ _02853_ _02858_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09088_ _03776_ _03777_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_169_Right_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output179_I net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08800__B2 as2650.stack\[14\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08039_ _02793_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11050_ as2650.stack\[0\]\[10\] _05461_ _05466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10001_ _04597_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10124__I _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07119__A1 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_150_Left_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08529__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_47_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10903_ _04778_ _05339_ _05340_ _05341_ _05342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_135_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10834_ _05275_ _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10426__A1 _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10794__I _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10765_ _05177_ _05222_ _05223_ _05225_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_54_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10696_ _05173_ _05181_ _05183_ _00812_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_129_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09044__A1 _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_147_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05605__A1 _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11317_ _00113_ clknet_leaf_105_wb_clk_i net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_50_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11248_ _00044_ clknet_leaf_135_wb_clk_i as2650.stack\[11\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08555__B1 _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09898__A3 _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11179_ _05547_ _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_120_1775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_87_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05740_ _00752_ net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_91_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07343__I _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05671_ _00665_ _00683_ _00684_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_114_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__B _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07410_ _02239_ _02240_ _02241_ _02094_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_72_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08390_ as2650.stack\[7\]\[14\] _02510_ _02513_ as2650.stack\[6\]\[14\] _03111_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ _02113_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08174__I _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ net68 net67 net69 _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_132_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07833__A2 _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_132_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05844__A1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09011_ _03702_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_132_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06223_ _01139_ _01140_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A1 _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06154_ _01125_ _01126_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold101 wbs_dat_i[18] net447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_125_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold112 wbs_dat_i[24] net458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_44_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06085_ net231 net250 _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09913_ _04554_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_1704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ as2650.trap as2650.irqs_latch\[4\] _04514_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_126_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09775_ _01887_ _02607_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06987_ _01898_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_1435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08726_ _03092_ _03424_ _03101_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05938_ _00745_ as2650.instruction_args_latch\[11\] _00941_ _00942_ _00943_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__08849__A1 as2650.stack\[11\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08313__A3 _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09510__A2 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08657_ as2650.stack\[8\]\[4\] _03302_ _03303_ as2650.stack\[9\]\[4\] _03130_ _03358_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05869_ _00862_ _00866_ net196 _00875_ net345 _00702_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_1_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07608_ _02390_ _02397_ _02398_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08588_ as2650.stack\[3\]\[2\] _03289_ _03290_ as2650.stack\[2\]\[2\] _03291_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10408__A1 _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07539_ wb_counter\[5\] _02342_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_27_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10550_ _05073_ _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_9_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09209_ _03881_ _03891_ _03894_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05835__A1 _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ as2650.stack\[2\]\[12\] _05039_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09577__A2 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__A4 _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11102_ _05445_ _05495_ _05500_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09329__A2 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_121_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11033_ as2650.stack\[0\]\[5\] _05451_ _05454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08001__A2 _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_138_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_138_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_19_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09501__A2 _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_169_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10817_ _05147_ _05258_ _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_83_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11797_ _00576_ clknet_leaf_28_wb_clk_i as2650.stack\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08208__B _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10748_ _04769_ _05142_ _05164_ _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_32_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05826__B2 as2650.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10029__I _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _04931_ _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_129_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09568__A2 _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput206 net206 la_data_out[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10178__A3 _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput217 net217 la_data_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08776__B1 _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput228 net228 last_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput239 net239 ram_enabled vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_107_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06242__I _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_15__f_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06910_ as2650.PC\[5\] _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07890_ as2650.indirect_target\[0\] _02635_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06003__A1 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09740__A2 _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ as2650.stack\[12\]\[1\] _01739_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06554__A2 _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _04242_ _04244_ _04245_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06772_ _01692_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_121_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_121_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10638__A1 _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08511_ _03197_ _03215_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05723_ _00735_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09491_ _01491_ _01021_ _04175_ _04176_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_78_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07503__A1 net165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08442_ _01276_ _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05654_ net239 _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_91_1689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _03070_ _03092_ _03094_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05585_ _00598_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11470__D _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07324_ net296 _02166_ _02160_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08833__S _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07255_ _02080_ _02103_ _02104_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06206_ _01117_ _01178_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_76_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09559__A2 _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07186_ _02048_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_76_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06137_ _01108_ _01109_ _00666_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_112_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input55_I ram_bus_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _01042_ _01049_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09827_ _02570_ _04502_ _04505_ _03534_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_96_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_1833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _02708_ _04439_ _04441_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_output211_I net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08709_ _03404_ _03405_ _03406_ _03407_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09689_ _04353_ _04374_ _03799_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09495__A1 _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11720_ _00504_ clknet_leaf_77_wb_clk_i as2650.regs\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05940__B _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11651_ _00435_ clknet_leaf_82_wb_clk_i as2650.regs\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09247__A1 _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08028__B _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11054__A1 _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ as2650.stack\[7\]\[3\] _05118_ _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11582_ _00366_ clknet_leaf_94_wb_clk_i as2650.regs\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10533_ _01685_ _01713_ _01970_ _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_68_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08542__I _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10464_ _04639_ _05026_ _05029_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10395_ _04736_ _04883_ _01423_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_1692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06784__A2 _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11016_ as2650.stack\[0\]\[0\] _05441_ _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_161_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08289__A2 _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11849_ net301 net168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09238__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_16_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11045__A1 _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09789__A2 _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_4_6__leaf_wb_clk_i clknet_leaf_35_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07040_ as2650.stack\[12\]\[13\] _01941_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07068__I _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09961__A2 _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08991_ _03682_ _03604_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_142_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07972__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06775__A2 _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ _02615_ _01765_ _02700_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08401__B _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07873_ _02634_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11465__D _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09612_ _04296_ _04297_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_108_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06824_ _01743_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_108_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09543_ _02565_ _04228_ _03726_ _03644_ _03774_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_116_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06755_ _01666_ _00727_ _01676_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_52_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05706_ _00718_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09474_ _04127_ _03928_ _04089_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_133_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06686_ _01353_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08425_ _03136_ _03139_ _03140_ _03144_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05637_ _00591_ _00643_ _00650_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_19_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08356_ net205 _01436_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_78_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07307_ net165 _02147_ _02148_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08287_ _03000_ _02617_ _03002_ net206 _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_85_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06463__A1 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07238_ _01561_ _02083_ _02085_ _02088_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_1691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07169_ net81 net114 _02036_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_output161_I net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _04749_ _04752_ _04755_ _04756_ _04758_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__08755__A3 _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07963__A1 _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_1718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_54_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11703_ _00487_ clknet_leaf_13_wb_clk_i as2650.stack\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08691__A2 _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11634_ _00418_ clknet_leaf_14_wb_clk_i as2650.stack\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11565_ _00349_ clknet_leaf_8_wb_clk_i as2650.stack\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09640__A1 _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09640__B2 _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06454__A1 _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10516_ as2650.stack\[1\]\[9\] _05060_ _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11496_ _00280_ clknet_leaf_136_wb_clk_i as2650.stack\[5\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10447_ _05017_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10002__A2 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10378_ _02893_ _01384_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_163_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_153_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_153_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06509__A2 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10042__I _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06540_ _00897_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10069__A2 _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07351__I _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06471_ _01198_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08210_ _01034_ _02948_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_116_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09190_ _00756_ _00874_ _00855_ _00717_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ as2650.indirect_target\[13\] _02757_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09631__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08072_ _01877_ _01862_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_128_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07023_ _01931_ _01756_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07945__A1 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08974_ _03626_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07526__I _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold16 _00124_ net360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_1505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ _02607_ _02683_ _02684_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold27 _00127_ net371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold38 _02395_ net382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold49 net450 net393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_58_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ as2650.insin\[3\] _02612_ _02620_ _01288_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_93_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input18_I bus_in_sid[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06807_ _01082_ _01573_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_155_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07787_ _02474_ _02554_ _02555_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_09526_ _03684_ _03680_ _03681_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06738_ _01658_ _01661_ _01527_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09457_ _04140_ _04142_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_109_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06669_ _01357_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_148_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08673__A2 _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11009__A1 _05391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08408_ _02666_ _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09388_ _04061_ _04063_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_4_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ _03060_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_43_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09622__A1 _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10232__A2 _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11350_ net383 clknet_leaf_107_wb_clk_i wb_counter\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10301_ _04164_ _04783_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11281_ _00077_ clknet_leaf_104_wb_clk_i net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_56_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10232_ _01460_ _01795_ _02585_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_56_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09925__A2 _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10163_ _04730_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10290__C _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ _04667_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08361__A1 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08267__I _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10996_ _05290_ as2650.regs\[4\]\[5\] _03104_ _05425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11727__CLK clknet_4_15__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09700__I2 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11617_ _00401_ clknet_leaf_120_wb_clk_i as2650.stack\[1\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09613__A1 _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11548_ _00332_ clknet_leaf_9_wb_clk_i as2650.stack\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11479_ _00263_ clknet_leaf_30_wb_clk_i as2650.debug_psu\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_0_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09916__A2 net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08730__I _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07774__C _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09047__B _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05971_ _00950_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_119_1809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07710_ _02473_ _02478_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_105_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08690_ _01830_ _03375_ _03389_ _03197_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_139_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08352__A1 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07641_ wb_counter\[25\] _02424_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_7_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07572_ _02358_ _02367_ net378 _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_50_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09311_ _03993_ _03996_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_152_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06523_ _01480_ _01482_ _01483_ _01293_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_76_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _03902_ _03906_ _03927_ _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06454_ _01387_ _01397_ _01416_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_139_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09173_ _03734_ _03854_ _03859_ _03733_ _03747_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_111_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06385_ _00862_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_146_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08124_ as2650.indirect_target\[11\] _01330_ _02848_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06418__A1 _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_135_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06969__A2 _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ as2650.ivectors_base\[2\] _02610_ _02809_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07006_ _01915_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_25_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_92_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09907__A2 net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10922__B1 _05359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07394__A2 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08957_ _03610_ _03616_ _03645_ _03648_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_07908_ _01546_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08888_ as2650.debug_psl\[0\] _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07192__S _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07839_ _00667_ _00677_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XANTENNA_output124_I net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10850_ _05290_ _00851_ _01525_ _04767_ _05291_ _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_49_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_49_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ net217 net216 net215 _01492_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_94_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10781_ as2650.stack\[6\]\[3\] _05232_ _05236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06657__A1 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11402_ _00186_ clknet_leaf_46_wb_clk_i as2650.indirect_target\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_62_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06335__I _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11333_ _00129_ clknet_leaf_154_wb_clk_i wb_counter\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_1458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11264_ _00060_ clknet_leaf_147_wb_clk_i net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__08550__I _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10215_ _04744_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_140_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11195_ as2650.stack\[9\]\[5\] _05557_ _05559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_145_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10146_ _04234_ _04236_ _04237_ _04238_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_78_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06593__B1 _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10077_ _04621_ _04668_ _04671_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08334__A1 _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10141__A1 _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10979_ _05396_ _05412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06170_ net56 _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_143_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08661__S _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05623__A2 _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09860_ _01737_ _04526_ _04529_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08811_ _03482_ _03505_ _03506_ _03103_ _02942_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09791_ _04439_ _04471_ _04472_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10380__A1 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05926__A3 _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08742_ _03434_ _03439_ _02549_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05954_ _00958_ _00646_ _00590_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_139_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07804__I _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08673_ _01830_ _03280_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10132__A1 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05885_ _00847_ _00890_ _00891_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08876__A2 _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07624_ _02407_ _02409_ _02411_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_85_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07555_ net394 _02344_ _02351_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08628__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09825__A1 _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06506_ _01467_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07486_ net83 _02060_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09225_ _03895_ _03899_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_98_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06437_ _01162_ _01365_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_40_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09156_ _02467_ _03648_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06368_ _01299_ _01301_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_161_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08107_ _02855_ _02857_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09087_ _01283_ _03592_ _03693_ _02920_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06299_ _01252_ _01256_ _01270_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08800__A2 _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08038_ _02633_ _02683_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_47_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_111_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08939__I0 _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10000_ _04595_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output241_I net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09989_ _01869_ _04603_ _04608_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10371__A1 _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05943__B _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07714__I _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10123__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06878__A1 _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10902_ _05275_ _05341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10833_ _05257_ _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09816__A1 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10764_ as2650.regs\[6\]\[5\] _05225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10977__A3 _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10695_ _05172_ _05181_ _05183_ _00884_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_clkbuf_leaf_150_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05605__A2 _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11316_ _00112_ clknet_leaf_102_wb_clk_i net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_1_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08280__I _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11247_ _00043_ clknet_leaf_136_wb_clk_i as2650.stack\[11\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_143_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11178_ _01713_ _01962_ _04522_ _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10362__A1 _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06949__B _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10129_ _04704_ _04705_ _04706_ _04707_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__06581__A3 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A1 _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08858__A2 _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10050__I _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05670_ _00669_ net50 _00670_ _00672_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_77_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__A2 _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07340_ _02162_ _02179_ _02180_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_161_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07294__A1 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07271_ _02118_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09010_ _01257_ _03701_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_132_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06222_ _01162_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_132_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold115_I wbs_dat_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07046__A1 _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06153_ as2650.insin\[3\] _01095_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold102 wbs_dat_i[14] net448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_160_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold113 wbs_dat_i[2] net459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_48_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11595__CLK clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06084_ _01063_ net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09912_ _04555_ _01637_ _04561_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_74_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09843_ _04517_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10353__A1 _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06986_ _01889_ _01897_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09774_ _02599_ _04455_ _04456_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05937_ _00744_ _00630_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08725_ _03091_ _03071_ _03090_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_119_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11056__I _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08849__A2 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08656_ as2650.stack\[11\]\[4\] _03308_ _03296_ as2650.stack\[10\]\[4\] _03357_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05868_ _00874_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09510__A3 _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07607_ net81 _02394_ _02385_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08587_ _01966_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05799_ _00662_ _00805_ _00808_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07538_ _02131_ _02336_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07285__A1 net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07469_ _02278_ wb_counter\[29\] _02272_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_92_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09208_ _00719_ _03892_ _01499_ _03893_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_169_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output191_I net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10480_ _05020_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output289_I net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07037__A1 _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09139_ as2650.debug_psl\[0\] _01780_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_121_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11101_ as2650.stack\[14\]\[2\] _05497_ _05500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11032_ _01834_ _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10344__A1 _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06488__C _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05771__A1 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06315__A3 _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_107_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_107_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_hold93_I wbs_dat_i[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10816_ _05255_ _05256_ _05257_ _05258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_11796_ _00575_ clknet_leaf_18_wb_clk_i as2650.stack\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11072__A2 _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10747_ _01584_ _01595_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10678_ _05173_ _05167_ _05170_ _00818_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_11_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07028__A1 _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07619__I _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput207 net207 la_data_out[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput218 net218 la_data_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput229 net229 last_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_107_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08878__C _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06003__A2 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06840_ _01759_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06771_ _01691_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_136_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05762__A1 _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08510_ _03198_ _03199_ _03214_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_121_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05722_ _00734_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09490_ _04036_ _04037_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_82_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08700__A1 _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08441_ _01727_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05653_ net59 _00666_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_118_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08372_ _02812_ _03093_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05584_ as2650.relative_cyc as2650.indirect_cyc _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_50_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07323_ _02136_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_119_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07254_ net277 _02095_ _02075_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_1586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10810__A2 _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09008__A2 _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06205_ net139 _01176_ _01177_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_144_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_1738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07185_ net89 net121 _02046_ _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_76_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06136_ _01104_ net52 _00671_ _00673_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_131_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06067_ _01040_ _01041_ _01044_ _00857_ _01047_ _01048_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_125_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08519__A1 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09744__I _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input48_I irqs[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10326__A1 _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ net181 _02480_ _04504_ _02483_ _02569_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07264__I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05753__A1 _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09757_ _04440_ _02640_ _03708_ _03710_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_5_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06969_ _01876_ _01881_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10629__A2 _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08708_ as2650.stack\[4\]\[6\] _02488_ _02495_ as2650.stack\[5\]\[6\] _02516_ _03407_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_154_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09688_ _03716_ _04366_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09495__A2 _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output204_I net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08639_ _03229_ _01792_ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_29_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11650_ _00434_ clknet_leaf_92_wb_clk_i as2650.regs\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _05080_ _05116_ _05121_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11581_ _00365_ clknet_leaf_92_wb_clk_i as2650.regs\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10532_ _01736_ _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10463_ as2650.stack\[2\]\[5\] _05027_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08758__A1 _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10394_ as2650.regs\[5\]\[6\] _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06233__A2 _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07430__A1 _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10317__A1 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11015_ _05440_ _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11290__CLK clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11848_ net301 net167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07249__A1 _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11779_ _00558_ clknet_leaf_4_wb_clk_i as2650.stack\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06472__A2 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_75_wb_clk_i clknet_4_15__leaf_wb_clk_i clknet_leaf_75_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08749__A1 _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_110_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__A1 _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08990_ _03600_ _03650_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07972__A2 _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07941_ _02606_ _01744_ _02699_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_62_1792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09174__A1 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ _01264_ _02633_ _01472_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__10503__I _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08921__A1 _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _01806_ _01559_ _03580_ _01568_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_108_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06823_ as2650.PC\[0\] as2650.PC\[1\] _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_108_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09542_ _03619_ _03671_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06754_ _01666_ _00935_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05705_ _00717_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_65_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07488__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06685_ _01599_ _01601_ _01613_ net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_09473_ _04144_ _04158_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_56_1596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05636_ _00591_ _00649_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08424_ as2650.stack\[15\]\[15\] _03141_ _03143_ as2650.stack\[14\]\[15\] _03117_
+ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_149_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08355_ _02606_ net205 _01438_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_24_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_78_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07306_ net134 _02149_ _02150_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08286_ _03013_ _03014_ _02622_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07237_ _02086_ net122 _02087_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07168_ _02038_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_1579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09401__A2 _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06119_ as2650.debug_psu\[5\] _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_105_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07099_ _01972_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_1578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output154_I net154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09809_ _04430_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05726__A1 _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08676__B1 _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11702_ _00486_ clknet_leaf_11_wb_clk_i as2650.stack\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06338__I _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06151__A1 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _00417_ clknet_leaf_114_wb_clk_i as2650.stack\[15\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08428__B1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11564_ _00348_ clknet_leaf_9_wb_clk_i as2650.stack\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10786__A1 _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09640__A2 _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06454__A2 _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10515_ _04645_ _05059_ _05061_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11495_ _00279_ clknet_leaf_127_wb_clk_i as2650.stack\[5\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold56_I net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10446_ _05016_ _04665_ _04622_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06206__A2 _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _01387_ _04792_ _04948_ _04950_ _04815_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_46_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_163_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06801__I _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07706__A2 _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08903__A1 _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10710__A1 _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_122_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_122_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07632__I _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ _01278_ _01152_ _01432_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_115_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08419__B1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08140_ as2650.ivectors_base\[9\] _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08463__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09631__A2 _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08071_ _02744_ _02823_ _02824_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_153_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07079__I _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07022_ as2650.debug_psu\[4\] _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_148_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07807__I _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08973_ _03631_ _03659_ _03660_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xhold17 net457 net361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_07924_ _02643_ _02682_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10233__I _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold28 wbs_dat_i[10] net372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold39 _00146_ net383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_97_1652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07855_ _02619_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06806_ _01131_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07786_ _01433_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06586__C _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09525_ _03683_ _03649_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_79_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06737_ _01543_ _01660_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08658__B1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08122__A2 _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06158__I _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09456_ _04115_ _04141_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06668_ _00180_ _01587_ _01597_ _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05619_ _00630_ _00632_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_08407_ _03127_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09387_ _04071_ _04072_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06599_ _01239_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_87_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05997__I _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ _01101_ _03059_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09622__A2 _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ as2650.instruction_args_latch\[8\] _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07633__A1 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10232__A3 _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08830__B1 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10300_ _01769_ _04774_ _04875_ _04876_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_132_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11280_ _00076_ clknet_leaf_103_wb_clk_i net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_61_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08189__A2 _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ _04358_ _04808_ _04793_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_56_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11193__A1 as2650.stack\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ _04733_ _04735_ _04738_ _04740_ _03658_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XTAP_TAPCELL_ROW_7_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_4_13__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10093_ _04643_ _04675_ _04680_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08548__I _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07452__I _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10995_ _04959_ _04960_ _05399_ _05424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_152_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07872__A1 _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_152_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11616_ _00400_ clknet_leaf_121_wb_clk_i as2650.stack\[1\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_169_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11547_ _00331_ clknet_leaf_8_wb_clk_i as2650.stack\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11478_ _00262_ clknet_leaf_31_wb_clk_i net181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10429_ _01382_ _04917_ _04999_ _05000_ _04756_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_81_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06531__I _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05938__A1 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11149__I _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10053__I _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05970_ _00747_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08886__C _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_105_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08352__A2 _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07640_ wb_counter\[23\] wb_counter\[24\] _02416_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_75_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07571_ net377 _02361_ _02368_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06522_ _01440_ _01303_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_117_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09310_ _03983_ _03994_ _03995_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_92_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06453_ _01404_ _01410_ _01412_ _01415_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_111_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09241_ _03910_ _03926_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_145_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_139_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09172_ _03857_ _03742_ _03743_ _03858_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_17_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06384_ _00899_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08123_ as2650.instruction_args_latch\[11\] _02740_ _02712_ _02873_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10228__I _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09080__A3 _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08054_ _01547_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07005_ as2650.PC\[11\] _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07537__I _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08040__A1 _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08956_ _03646_ _03647_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input30_I bus_in_timers[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07907_ _01427_ _02664_ _02665_ _02667_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_08887_ _03102_ _03560_ _03579_ _03534_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_58_1422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07838_ _02449_ _02605_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_1499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output117_I net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07769_ as2650.stack\[12\]\[13\] _02534_ _02537_ as2650.stack\[13\]\[13\] _02538_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_49_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09508_ _00833_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_91_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10780_ _05080_ _05230_ _05235_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10989__A1 _05347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09439_ _04108_ _04124_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_140_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06616__I _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11401_ _00185_ clknet_leaf_46_wb_clk_i as2650.indirect_target\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_145_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08803__B1 _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05617__B1 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11332_ _00128_ clknet_leaf_147_wb_clk_i as2650.wb_hidden_rom_enable vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_127_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11263_ _00059_ clknet_leaf_134_wb_clk_i net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__11166__A1 as2650.stack\[13\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08031__A1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10214_ _04711_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11194_ _05449_ _05556_ _05558_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_145_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10913__A1 _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10145_ _04723_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06593__A1 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06593__B2 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10076_ as2650.stack\[3\]\[0\] _04670_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07182__I _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10978_ _05296_ _05409_ _05410_ _05411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09598__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09837__I _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06820__A2 _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11157__A1 _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10904__A1 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_1582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08810_ _03009_ _03096_ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09770__A1 _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09790_ _01316_ _04429_ _04465_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_139_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ _03435_ _03436_ _03437_ _03438_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_119_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05953_ as2650.page_reg\[0\] _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09522__A1 _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08672_ _03193_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05884_ _00845_ as2650.regs\[6\]\[2\] _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07623_ net85 _02410_ _02401_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08089__A1 _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ wb_counter\[8\] _02354_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06505_ _01290_ _01466_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_158_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07485_ _01561_ _02059_ _02302_ _02063_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_9_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _03907_ _03908_ _03909_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_98_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06436_ _01348_ _01375_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_57_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06367_ _01250_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09155_ _01167_ _02564_ _03841_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_66_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08106_ _02856_ _02829_ _02838_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_146_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06298_ _01259_ _01261_ _01269_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09086_ _03775_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08037_ _02791_ _02661_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08939__I1 _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09988_ as2650.stack\[4\]\[7\] _04604_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output234_I net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08939_ _00686_ _01357_ _01210_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_150_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06120__B _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10901_ _04174_ _04963_ _05340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_64_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10832_ _05264_ _04964_ _05269_ _05273_ _05274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_67_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10763_ _05174_ _05222_ _05223_ _05224_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_95_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10694_ _05171_ _05181_ _05183_ _00860_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_118_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07886__B _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_147_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11315_ _00111_ clknet_leaf_140_wb_clk_i net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_73_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_147_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05605__A3 _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11246_ _00042_ clknet_leaf_135_wb_clk_i as2650.stack\[11\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08555__A2 _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09752__A1 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11177_ _05477_ _05541_ _05546_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_1777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10128_ as2650.cycle\[10\] _01695_ _01528_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_78_1639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10059_ as2650.stack\[10\]\[12\] _04657_ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06318__A1 _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10114__A2 _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_29_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_82_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09060__C _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07270_ _02117_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07294__A2 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08491__A1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06221_ _01191_ _01193_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_2_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09035__A3 _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06152_ _01117_ _01124_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_91_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold108_I wbs_dat_i[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07046__A2 _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08471__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08243__B2 net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold103 wbs_dat_i[19] net449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold114 wbs_adr_i[21] net460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_06083_ net350 _00930_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _04556_ net150 _04557_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09842_ net46 as2650.irqs_latch\[3\] _04514_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09773_ _01887_ _02599_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06985_ _01843_ _01894_ _01896_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_119_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08724_ _03065_ _03400_ _03402_ _03422_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05936_ _00940_ _00627_ _00629_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08655_ _03352_ _03353_ _03354_ _03355_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05867_ _00873_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07606_ wb_counter\[18\] _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_49_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08586_ _01690_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05798_ _00743_ as2650.instruction_args_latch\[5\] _00806_ _00807_ _00808_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_152_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07537_ _02340_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08482__A1 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07285__A2 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07468_ net110 _02279_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09207_ _01493_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06419_ _01345_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07399_ _02124_ _01887_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07198__S _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09138_ _03661_ _03659_ _03660_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08381__I _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output184_I net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08785__A2 _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09069_ _01755_ _02608_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_163_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11100_ _05443_ _05495_ _05499_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11031_ _05449_ _05450_ _05452_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10344__A2 _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05771__A2 as2650.instruction_args_latch\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06315__A4 _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06720__A1 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10815_ _01750_ _03725_ _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_83_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11795_ _00574_ clknet_leaf_5_wb_clk_i as2650.stack\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold86_I wbs_dat_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _05112_ _05208_ _05213_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08473__A1 _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09670__B1 _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_147_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_147_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _04904_ _05173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_168_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08225__A1 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06804__I _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09973__A1 _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A2 _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 net208 la_data_out[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput219 net219 la_data_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_1390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06787__A1 _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10583__A2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_166_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09725__A1 _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11229_ _00025_ clknet_leaf_133_wb_clk_i as2650.stack\[12\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_125_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10061__I _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06770_ _01690_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05721_ net345 _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08161__B1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08700__A2 _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08440_ _03156_ _03157_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05652_ _00665_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_59_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05583_ _00594_ _00596_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_08371_ net212 _01439_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ _02155_ wb_counter\[8\] _02164_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08464__A1 as2650.ivectors_base\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_119_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07253_ _02082_ _02100_ _02102_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06204_ net62 _01080_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06714__I _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07184_ _02047_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06135_ _01104_ _01105_ _01106_ _01107_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_147_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06066_ _01041_ _00836_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09716__A1 _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09825_ _01838_ _02485_ _04503_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09756_ _01872_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_154_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06968_ _01787_ _01878_ _01880_ _01842_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08707_ as2650.stack\[7\]\[6\] _01688_ _01964_ as2650.stack\[6\]\[6\] _03406_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05919_ _00911_ _00915_ _00919_ _00923_ _00734_ _00703_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_09687_ _04372_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_119_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06899_ _01815_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_94_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _01788_ _02464_ _03339_ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06702__A1 net241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07280__I _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08569_ _01744_ _03243_ _03268_ _02557_ _03272_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_166_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10600_ as2650.stack\[7\]\[2\] _05118_ _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07258__A2 _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08455__A1 _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11580_ _00364_ clknet_leaf_94_wb_clk_i as2650.regs\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10531_ _04663_ _05065_ _05070_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10462_ _04635_ _05026_ _05028_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09000__I _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__A2 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10393_ _04939_ _04787_ _04961_ _04724_ _04966_ _04771_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__09935__I _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07430__A2 _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09183__A2 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11014_ _05437_ _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_99_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11435__CLK clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08930__A2 _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07497__A2 _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_1654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11847_ net301 net166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07249__A2 net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11778_ _00557_ clknet_leaf_3_wb_clk_i as2650.stack\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10729_ as2650.stack\[8\]\[8\] _05203_ _05204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06472__A3 _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09946__A1 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A2 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10056__I _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__A2 _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07940_ _01719_ _02645_ _02681_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09066__B _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_1801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_44_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_44_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09174__A2 _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ _01319_ _01325_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09610_ _01754_ as2650.debug_psl\[2\] _03732_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08921__A2 _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06822_ _01724_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_108_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09541_ _03672_ _03639_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_69_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06753_ net246 _01007_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05704_ _00716_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07488__A2 _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09472_ _04143_ _04128_ _04131_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06684_ _01551_ _01610_ _01611_ _01612_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_133_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08685__A1 _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08423_ _03142_ _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05635_ _00644_ _00647_ _00648_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ _02714_ _03075_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10244__A1 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ _02121_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08285_ _03007_ _02846_ _01256_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06999__A1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07236_ _02011_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06463__A3 _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05671__A1 _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09937__A1 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07167_ net80 net113 _02036_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input60_I rom_bus_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10547__A2 _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06118_ net44 net43 net46 net45 _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_100_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07098_ _01928_ _01986_ _01991_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_112_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06049_ wb_reset_override_en net33 _01032_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_1_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09165__A2 _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output147_I net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09808_ net214 _04449_ _04488_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i clknet_4_15__leaf_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09739_ _04403_ _04423_ _04372_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11701_ _00485_ clknet_leaf_11_wb_clk_i as2650.stack\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06151__A2 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11632_ _00416_ clknet_leaf_114_wb_clk_i as2650.stack\[15\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08428__A1 _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10235__A1 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11563_ _00347_ clknet_leaf_8_wb_clk_i as2650.stack\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08055__B _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06354__I _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10514_ as2650.stack\[1\]\[8\] _05060_ _05061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_150_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11494_ _00278_ clknet_leaf_39_wb_clk_i as2650.stack\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_96_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10445_ _01712_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10538__A2 _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10376_ _04949_ _04729_ _04792_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_103_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10604__I _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07706__A3 _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08903__A2 _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07913__I _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10710__A2 _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09703__I1 net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06529__I _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08667__A1 _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_116_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10226__A1 _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09092__A1 _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ as2650.ivectors_base\[3\] _02610_ _02809_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05653__A1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07021_ _01715_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10529__A2 _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08412__C _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08972_ _03635_ _03662_ _03663_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_45_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07923_ _02642_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold18 net99 net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold29 net73 net373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_157_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07854_ _01124_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06805_ _01721_ _01725_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_135_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07785_ _01172_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_135_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09524_ _03594_ _03842_ _04209_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06736_ _01606_ _00805_ _01659_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_17_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09455_ _04117_ _04119_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_52_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06667_ _01593_ _01594_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08406_ _03105_ _03122_ _03126_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05618_ _00631_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_30_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_130_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09386_ _04048_ _04064_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06598_ _01544_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_35_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08337_ _03058_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08268_ _01480_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ net161 net94 _02069_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08199_ _02933_ _02934_ _02936_ _02940_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10230_ _04709_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_56_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08594__B1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10161_ _04739_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_63_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05947__A2 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_4_0__f_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10092_ as2650.stack\[3\]\[7\] _04676_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_143_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07733__I _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06349__I as2650.cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08649__A1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08649__B2 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10994_ _05408_ _05422_ _05423_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10456__A1 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A1 _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11615_ _00399_ clknet_leaf_121_wb_clk_i as2650.stack\[1\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_169_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11546_ _00330_ clknet_leaf_9_wb_clk_i as2650.stack\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05635__A1 _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11477_ _00261_ clknet_leaf_30_wb_clk_i as2650.debug_psu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _03783_ _04861_ _04917_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_164_Right_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11184__A2 _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10359_ _04933_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05938__A2 as2650.instruction_args_latch\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08352__A3 _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ _02292_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06521_ _01446_ _01481_ _01294_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07312__A1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10998__A2 _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _03912_ _03925_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06452_ _01413_ _01414_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__08474__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09171_ _01389_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06383_ _00834_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09065__B2 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08122_ as2650.indirect_target\[11\] _02680_ _02844_ _02871_ _02872_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_135_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08812__A1 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_135_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08053_ as2650.indirect_target\[6\] _02654_ _02657_ _02792_ _02807_ _02808_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_43_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07004_ _01871_ _01913_ _01914_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06426__I0 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10922__A2 _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08955_ _03609_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_102_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07906_ _02666_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08886_ _03277_ _03577_ _03578_ _03101_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_97_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input23_I bus_in_sid[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07837_ as2650.insin\[0\] _02596_ _02600_ _02603_ _02604_ _02605_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_100_1594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07551__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07768_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09507_ _01856_ _04186_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06719_ _01639_ _01644_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _02467_ _01198_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_66_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09438_ _04120_ _04123_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08384__I _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05865__A1 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09369_ _04047_ _04053_ _04054_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XANTENNA__09056__A1 _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11400_ _00184_ clknet_leaf_47_wb_clk_i as2650.indirect_target\[4\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_1_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08803__A1 _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11331_ net371 clknet_leaf_145_wb_clk_i net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_132_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07728__I _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A2 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11262_ _00058_ clknet_leaf_148_wb_clk_i net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__06632__I _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10213_ _04757_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11193_ as2650.stack\[9\]\[4\] _05557_ _05558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_145_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_120_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10144_ _04695_ _04700_ _04722_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_TAPCELL_ROW_145_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06593__A2 _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10075_ _04669_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_141_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07542__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10429__A1 _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10977_ _03813_ as2650.regs\[4\]\[1\] _03104_ _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_15_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09047__A1 _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09598__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__I0 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05608__A1 as2650.indirect_target\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05608__B2 as2650.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10601__A1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11529_ _00313_ clknet_leaf_72_wb_clk_i net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_41_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_130_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10064__I _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08740_ as2650.stack\[15\]\[7\] _03428_ _03429_ as2650.stack\[14\]\[7\] _02517_ _03438_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05952_ _00645_ as2650.extend as2650.instruction_args_latch\[13\] _00957_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08671_ _03348_ _03369_ _03371_ _03103_ _02942_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05883_ as2650.regs\[2\]\[2\] _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10132__A3 _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ _02339_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07553_ _02353_ _02349_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__A2 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06504_ _01465_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07484_ net72 _02060_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09223_ _03887_ _03889_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_1742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06435_ _01162_ _01338_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_107_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09038__A1 _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09154_ _01152_ _01195_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_17_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06366_ _01316_ _01329_ _01330_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ _02826_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08797__B1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09085_ _03774_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_32_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06297_ _01265_ _01268_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08036_ _02790_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput90 net422 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08549__B1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ _01853_ _04603_ _04607_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08938_ _00662_ _01373_ _01225_ _03629_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_99_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07283__I _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10659__A1 _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output227_I net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10659__B2 _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08869_ _01934_ _03535_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__06327__A2 _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__A1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10900_ _05336_ _05337_ _05338_ _05339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08721__B1 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ as2650.chirpchar\[0\] _05271_ _05272_ _05273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10762_ as2650.regs\[6\]\[4\] _05224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06627__I _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10693_ _05163_ _05181_ _05183_ _00842_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_47_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06263__A1 _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11314_ _00110_ clknet_leaf_102_wb_clk_i net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05605__A4 _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11245_ _00041_ clknet_leaf_136_wb_clk_i as2650.stack\[11\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_1555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10898__A1 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11176_ as2650.stack\[13\]\[15\] _05542_ _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10127_ _01695_ _04373_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_101_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_1789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09504__A2 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _04626_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06318__A2 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07515__A1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_69_wb_clk_i clknet_4_13__leaf_wb_clk_i clknet_leaf_69_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05829__A1 _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_1758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06220_ _01192_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08779__B1 _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06151_ _01122_ _01123_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_93_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08243__A2 _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold104 wbs_dat_i[8] net450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_79_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06272__I _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold115 wbs_dat_i[0] net461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_06082_ _01051_ _01056_ _01058_ _01061_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_123_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09910_ _04555_ _01626_ _04560_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_1509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09841_ _02693_ _00010_ _04516_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09743__A2 _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10522__I _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ net199 _04449_ _04454_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06984_ _01895_ _01849_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _03403_ _03420_ _03421_ _03374_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05935_ _00625_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_87_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ as2650.stack\[4\]\[4\] _03302_ _03303_ as2650.stack\[5\]\[4\] _02519_ _03355_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05866_ _00872_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_68_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07605_ wb_counter\[17\] _02392_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08585_ _01443_ _03057_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05797_ _00743_ _00780_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08148__B _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07536_ _02339_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10813__A1 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07467_ _02277_ _02288_ _02289_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_162_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09206_ _00755_ _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06418_ _00738_ _01340_ _01342_ _01363_ _01381_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_17_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07398_ net114 _02149_ _02213_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09137_ _03610_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06349_ as2650.cycle\[6\] _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_103_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06245__A1 _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09068_ _03403_ _03756_ _03758_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output177_I net177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07993__A1 _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _02683_ _02774_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11030_ as2650.stack\[0\]\[4\] _05451_ _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06910__I as2650.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__A2 _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08170__A1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07741__I _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10814_ _01579_ _01750_ _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_28_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11794_ _00573_ clknet_leaf_5_wb_clk_i as2650.stack\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10745_ as2650.stack\[8\]\[15\] _05209_ _05213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09670__A1 _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08473__A2 _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09670__B2 _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10676_ _05172_ _05167_ _05170_ _00890_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09973__A2 _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput209 net209 la_data_out[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_65_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07984__A1 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_116_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_116_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_112_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07916__I _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11228_ _00024_ clknet_leaf_16_wb_clk_i as2650.stack\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11159_ _05523_ _05536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_159_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05720_ _00699_ _00667_ _00677_ _00732_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_121_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_121_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05651_ as2650.wb_hidden_rom_enable as2650.cpu_hidden_rom_enable _00665_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_37_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11048__A1 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03071_ _03090_ _03091_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_19_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06267__I _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05582_ _00595_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_54_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07321_ _01119_ _02147_ _02148_ _02163_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold120_I wbs_stb_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07252_ _02090_ _02101_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06203_ net42 _01154_ _01175_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08216__A2 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07183_ net88 net120 _02046_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09413__A1 _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06134_ net40 _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07975__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05825__I1 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06065_ _01045_ _01046_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09716__A2 _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09824_ _03755_ _03120_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i clknet_4_14__leaf_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06967_ _01879_ _01793_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09755_ _02588_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08706_ as2650.stack\[0\]\[6\] _02488_ _02495_ as2650.stack\[1\]\[6\] _02502_ _03405_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05918_ _00922_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09686_ as2650.cycle\[8\] _01539_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_119_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06898_ _01812_ _01814_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_154_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07561__I _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08637_ _01792_ _03243_ _03338_ _03242_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_55_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05849_ _00844_ _00846_ net195 _00856_ net346 _00703_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XTAP_TAPCELL_ROW_29_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08568_ _01444_ _03270_ _03271_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_49_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ _02321_ _02325_ _02326_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09652__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08499_ _02517_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10530_ as2650.stack\[1\]\[15\] _05066_ _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_86_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10461_ as2650.stack\[2\]\[4\] _05027_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09404__A1 _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _04159_ _04779_ _04965_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_81_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06640__I _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11013_ _05438_ _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_161_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__A1 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11777_ _00556_ clknet_leaf_3_wb_clk_i as2650.stack\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06457__A1 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10728_ _05190_ _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10659_ _04961_ _05156_ _05157_ _04966_ _05158_ _05160_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_TAPCELL_ROW_114_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06472__A4 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06209__A1 _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_110_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_110_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11168__I _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07870_ _01334_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08382__B2 _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ _01725_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_108_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06932__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ _01199_ _03831_ _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06752_ _00738_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_69_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08134__B2 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05703_ as2650.regs\[1\]\[7\] as2650.regs\[5\]\[7\] _00715_ _00716_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_13_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_13_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09471_ _04144_ _04152_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06683_ _01530_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_149_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08422_ _01966_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06696__A1 net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05634_ as2650.instruction_args_latch\[15\] _00647_ _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_153_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_120_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08353_ net206 _01436_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_24_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_24_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09634__A1 _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07304_ _02118_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08284_ _02997_ _03012_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_60_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ net67 _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_61_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ _02037_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07948__A1 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06117_ net48 net47 net49 _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_48_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_1813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07097_ as2650.stack\[11\]\[11\] _01987_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input53_I ram_bus_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06620__A1 _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ wb_reset_override wb_reset_override_en _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_58_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09570__B1 _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ _02484_ _04487_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07999_ _02748_ _02001_ _02755_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_96_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_2_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09738_ _04408_ _04422_ _04368_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09669_ _04353_ _04354_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08676__A2 _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11700_ _00484_ clknet_leaf_10_wb_clk_i as2650.stack\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10483__A2 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11631_ _00415_ clknet_leaf_114_wb_clk_i as2650.stack\[15\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09625__A1 _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08428__A2 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11562_ _00346_ clknet_leaf_9_wb_clk_i as2650.stack\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10513_ _05047_ _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11493_ _00277_ clknet_leaf_39_wb_clk_i as2650.stack\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_150_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05662__A2 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10444_ _04990_ _04787_ _05011_ _04724_ _05015_ _04771_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_61_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_139_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10375_ _04216_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_103_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08071__B _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06370__I _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06611__A1 net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_148_Left_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09703__I2 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09864__A1 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08419__A2 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09616__A1 _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_116_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06545__I _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10067__I _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_131_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_131_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_157_Left_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07020_ _01871_ _01928_ _01929_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09856__I _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09919__A2 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07376__I _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06280__I _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ _01557_ _01779_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07922_ _02646_ _02681_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold19 _02313_ net363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_100_1710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08355__A1 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09552__B1 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ _02611_ _02618_ _02004_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10162__B2 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_166_Left_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06804_ _01724_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07784_ _02523_ _02544_ _02552_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06735_ _01640_ _01026_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09523_ _01200_ _04202_ _04203_ _04208_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_116_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08658__A2 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09454_ _04135_ _04139_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06666_ _01596_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_137_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05617_ as2650.indirect_target\[12\] _00626_ _00628_ as2650.PC\[12\] _00631_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08405_ _03123_ _03125_ _03102_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09385_ _04051_ _04052_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06597_ _01543_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_164_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_47_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08336_ _03057_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08267_ _02933_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_43_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08830__A2 _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07218_ _02071_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08198_ _02937_ _02939_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08969__I0 _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _02027_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_56_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10160_ _01237_ _01099_ _04186_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_105_1643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10091_ _04641_ _04675_ _04679_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_7_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08346__A1 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09543__B1 _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10993_ _05359_ _05412_ _05416_ as2650.regs\[0\]\[4\] _05423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_156_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07321__A2 _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06380__I0 _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08066__B _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07872__A3 _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_152_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11614_ _00398_ clknet_leaf_124_wb_clk_i as2650.stack\[1\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08282__B1 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11545_ _00329_ clknet_leaf_117_wb_clk_i as2650.stack\[4\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11476_ _00260_ clknet_leaf_28_wb_clk_i as2650.debug_psu\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _01664_ _04848_ _04997_ _04998_ _04729_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10615__I _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_1444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10358_ _04772_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09625__B _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10289_ _02894_ _01406_ _01408_ _04865_ _04754_ _04866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_40_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10144__A1 _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_66_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06520_ _01233_ _01273_ _01287_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07312__A2 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06451_ _01411_ _01365_ _01366_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09170_ _03856_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_139_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06382_ _00924_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09065__A2 _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08121_ _02867_ _02870_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07076__A1 _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08273__B1 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08052_ _02698_ _02806_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07003_ as2650.stack\[12\]\[10\] _01884_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07379__A2 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06426__I1 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10383__A1 _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08954_ _03605_ _03606_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07834__I _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07905_ _01304_ _01483_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10135__A1 _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08885_ _02656_ _03240_ _03343_ _01936_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_07836_ _02462_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_input16_I bus_in_serial_ports[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07767_ _02535_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09506_ as2650.debug_psl\[6\] _02477_ _04191_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06718_ _01604_ _01643_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_49_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07698_ _01281_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_94_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09437_ _04121_ _04122_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06649_ _01585_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09368_ _04012_ _04016_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08319_ _03029_ _03042_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09299_ _03871_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_62_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11330_ net407 clknet_leaf_147_wb_clk_i wb_io3_test vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06814__A1 _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11261_ _00057_ clknet_leaf_149_wb_clk_i net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10212_ _01415_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11192_ _05550_ _05557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10374__A1 _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10143_ _04698_ _04721_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_145_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07744__I _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10074_ _04666_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_141_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10126__A1 _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09819__B2 _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10429__A2 _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09295__A2 _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10976_ _05403_ _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07058__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09598__A3 _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06805__A1 _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11528_ _00312_ clknet_leaf_73_wb_clk_i net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_164_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11459_ _00243_ clknet_leaf_42_wb_clk_i as2650.PC\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I bus_in_gpios[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05951_ _00747_ _00939_ _00955_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_4
XANTENNA__10117__A1 _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05792__A1 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ _03086_ _03370_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05882_ _00888_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08686__S _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05919__I0 _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07621_ wb_counter\[21\] _02408_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07552_ wb_counter\[7\] _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_85_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08485__I _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06503_ _01464_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07483_ _02237_ net427 _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06434_ _01388_ _01340_ _01342_ _01394_ _01396_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09222_ _03887_ _03889_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_98_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09038__A2 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_98_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09153_ _02469_ _03839_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_40_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06365_ _01254_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_133_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08104_ _02839_ _02854_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06733__I _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09084_ _01197_ _01230_ _03772_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_114_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08797__B2 as2650.stack\[9\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06296_ _01267_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08035_ _02789_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_86_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput80 net380 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput91 net415 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09986_ as2650.stack\[4\]\[6\] _04604_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08937_ _01607_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_102_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08868_ _02748_ _02882_ _03053_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_118_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08721__A1 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08721__B2 _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output122_I net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07819_ _02580_ _02561_ _02587_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_54_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ _02508_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_169_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10830_ _04777_ _05272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10761_ _05216_ _05223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_94_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10692_ _05182_ _05183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09029__A2 _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07739__I _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08788__A1 _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07460__A1 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ _00109_ clknet_leaf_102_wb_clk_i net280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11244_ _00040_ clknet_leaf_39_wb_clk_i as2650.stack\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10347__A1 _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11175_ _05475_ _05541_ _05545_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10126_ _01478_ _01503_ _03715_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_98_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10114__B _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _04624_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06318__A3 _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06818__I _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_80_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10959_ _05261_ _05393_ _05394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10822__A2 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_132_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06150_ net61 _01111_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_81_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_38_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_38_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_147_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10075__I _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ net230 _01060_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xhold105 wbs_dat_i[26] net451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold116 wbs_dat_i[17] net462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10338__B2 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09840_ net45 _00010_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10803__I _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08400__B1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i clknet_4_13__leaf_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09771_ _02473_ _04453_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06983_ _01890_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_33_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ _01848_ _02595_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05934_ _00938_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_119_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08653_ as2650.stack\[7\]\[4\] _03308_ _03296_ as2650.stack\[6\]\[4\] _03354_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05865_ _00715_ as2650.regs\[4\]\[1\] _00871_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__10510__A1 as2650.stack\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07604_ _02390_ _02393_ net382 _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05796_ _00779_ _00617_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08584_ _03284_ _03285_ _03286_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_117_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07535_ _02319_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_152_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07466_ net286 _02282_ _02275_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06417_ _01367_ _01380_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09205_ _00757_ _01499_ _01494_ _00718_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07397_ _02220_ _02229_ _02230_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08164__B _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06348_ _01313_ _01248_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09136_ _03822_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06245__A2 _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07442__A1 net282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09067_ _01755_ _03757_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06279_ _01250_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_103_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05599__A4 _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08018_ _02770_ _01829_ _02773_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__07993__A2 _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10329__A1 _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _04595_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10501__A1 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08170__A2 _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11862_ net173 net264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09014__I _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10813_ _01697_ _04300_ _05255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_0_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11793_ _00572_ clknet_leaf_19_wb_clk_i as2650.stack\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10744_ _05110_ _05208_ _05212_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__A2 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10675_ _04874_ _05172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06236__A2 _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08630__B1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05995__A1 net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11227_ _00023_ clknet_leaf_39_wb_clk_i as2650.stack\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05717__I _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11158_ _05521_ _05535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_125_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10109_ _04659_ _04687_ _04690_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11089_ _05178_ _05487_ _05488_ _05491_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_95_1730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_121_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_159_Right_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08161__A2 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05650_ _00663_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_110_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05581_ as2650.cycle\[0\] as2650.cycle\[4\] as2650.cycle\[6\] _00595_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_07320_ net136 _02149_ _02150_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07251_ wb_counter\[1\] _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_119_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06202_ _01174_ _01133_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07182_ _02035_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold113_I wbs_dat_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10559__A1 _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06133_ _00673_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_147_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11220__A2 _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09594__I _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07975__A2 _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06064_ as2650.indirect_target\[0\] _00635_ _00594_ as2650.cycle\[4\] _01046_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_112_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09177__A1 _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05627__I _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09823_ net306 _02791_ _04501_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09754_ _04431_ _04437_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06966_ _01877_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_119_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08705_ as2650.stack\[3\]\[6\] _01688_ _01964_ as2650.stack\[2\]\[6\] _03404_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_94_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05917_ _00690_ as2650.regs\[4\]\[4\] _00921_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09685_ _04363_ _04367_ _04368_ _04370_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_96_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06897_ _00602_ _01790_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08636_ _03324_ _03335_ _03336_ _03337_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05848_ _00855_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_139_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08567_ _01720_ _01762_ _01128_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05779_ as2650.regs\[1\]\[5\] as2650.regs\[5\]\[5\] _00789_ _00790_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09101__A1 _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07518_ net83 _02323_ _02293_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ as2650.stack\[7\]\[0\] _02508_ _02540_ as2650.stack\[6\]\[0\] _03203_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09652__A2 _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07663__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08606__C _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_21_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07449_ _02187_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10708__I _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _05020_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output287_I net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07415__A1 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09119_ _03159_ _02739_ _03708_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10391_ _01823_ _04932_ _04962_ _04964_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_143_1510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_1630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05977__A1 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08915__A1 _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07718__A2 _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ _05437_ _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10722__A1 _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07752__I _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold91_I _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11776_ _00555_ clknet_leaf_116_wb_clk_i as2650.stack\[14\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09643__A2 _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07654__A1 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10727_ _05188_ _05202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08851__B1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10658_ as2650.regs\[1\]\[5\] _05160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_114_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06209__A2 _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10589_ as2650.stack\[15\]\[15\] _05106_ _05113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_110_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08906__A1 _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06820_ _01716_ _01737_ _01740_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06393__A1 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06751_ _01664_ _01627_ _01672_ _01673_ net172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_69_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08134__A2 _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05702_ as2650.debug_psl\[4\] _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_91_1435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06682_ _01050_ _01551_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06278__I _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09470_ _04144_ _04152_ _04155_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_56_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08421_ _01691_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_153_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05633_ _00646_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_133_1745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07893__A1 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_53_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08352_ net207 _02619_ _01439_ _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_110_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09634__A2 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_24_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07303_ _02112_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_11_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08283_ _02998_ _02637_ _03009_ _03010_ _03011_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07234_ _02084_ net159 _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ net79 net106 _02036_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06116_ as2650.cycle\[11\] _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06741__I _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07096_ _01913_ _01986_ _01990_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06047_ _01031_ net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06620__A2 _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input46_I irqs[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09570__A1 _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09806_ _02552_ _04464_ _04486_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09570__B2 _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _02638_ _02752_ _02754_ _01320_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_57_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09737_ _04419_ _04421_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_2_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06949_ _01844_ _01827_ _01860_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11094__I _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09668_ _01749_ _01191_ _01342_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_167_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08619_ _03076_ _03082_ _03084_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_output202_I net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09599_ _04282_ _03731_ _04283_ _04284_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08617__B _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11630_ _00414_ clknet_leaf_126_wb_clk_i as2650.stack\[15\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07636__A1 wb_counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11561_ _00345_ clknet_leaf_89_wb_clk_i as2650.stack\[10\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10512_ _05045_ _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11492_ _00276_ clknet_leaf_15_wb_clk_i as2650.stack\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10443_ _05013_ _05014_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05662__A3 _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11196__A1 _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08061__A1 _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10374_ _01648_ _04793_ _04946_ _04947_ _04811_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_163_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09561__A1 _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11120__A1 _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06678__A2 _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07431__B _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09202__I _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07627__A1 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08824__B1 _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11759_ _00538_ clknet_leaf_99_wb_clk_i as2650.regs\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06602__A2 _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08970_ _03659_ _03660_ _03661_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xclkbuf_leaf_100_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_100_wb_clk_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07921_ _00678_ _01743_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_157_1509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08355__A2 net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07852_ as2650.insin\[2\] _02612_ _02617_ _01288_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__06366__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06803_ _01722_ _01723_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput1 bus_in_gpios[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07783_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09304__A1 _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09522_ _01168_ _04204_ _04207_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06734_ net244 _01007_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06118__A1 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07866__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09453_ _04138_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_133_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06665_ _01590_ _01594_ _01592_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08404_ _02927_ _03124_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05616_ _00625_ _00627_ _00629_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09384_ _04057_ _04068_ _04069_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_06596_ _01005_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08335_ _01131_ _02554_ _02555_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_129_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08266_ _02974_ _02996_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_144_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07217_ net160 net83 _02069_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08197_ _01316_ _02938_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06471__I _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07148_ net103 net137 _02025_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_56_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10925__A1 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07079_ _01972_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output152_I net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10090_ as2650.stack\[3\]\[6\] _04676_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09543__A1 _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08346__A2 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10153__A2 _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07157__I0 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _05349_ _05409_ _05421_ _05422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06380__I1 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11613_ _00397_ clknet_leaf_129_wb_clk_i as2650.stack\[1\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_152_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11544_ _00328_ clknet_leaf_118_wb_clk_i as2650.stack\[4\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11475_ _00259_ clknet_leaf_29_wb_clk_i as2650.debug_psu\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_hold54_I net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ _04279_ _04806_ _04858_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_123_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10357_ _04773_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_143_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10288_ _02893_ _02905_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_109_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09625__C _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08101__I _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07148__I0 net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09298__B1 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06450_ _01358_ _01374_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__A1 _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06381_ _01345_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_139_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08120_ _02789_ _01908_ _02869_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09867__I _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08051_ _02736_ _01456_ _02805_ _02724_ as2650.indirect_target\[6\] _02806_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_86_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07002_ _01912_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10907__A1 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__A2 _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09773__A1 _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06426__I2 net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06587__A1 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08953_ _03622_ _03639_ _03643_ _03644_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07904_ _01576_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08884_ _03561_ _03576_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06339__A1 _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07835_ _02602_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07000__A2 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_16_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_155_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07139__I0 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07766_ _02497_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09828__A2 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07850__I _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06894__C _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ _04189_ _04190_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06717_ _01642_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07839__A1 _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07697_ _02465_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09436_ _03915_ _04106_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06466__I _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06648_ _01239_ _01584_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_109_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09367_ _04048_ _04051_ _04052_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_06579_ _01196_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_35_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08318_ _02935_ _02937_ _02905_ _01449_ _03041_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__08264__A1 _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09298_ _01013_ _00898_ _00875_ _00913_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_69_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_25_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08249_ _02974_ _02982_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11260_ _00056_ clknet_leaf_148_wb_clk_i net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_10211_ _04786_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ _05548_ _05556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10142_ _04714_ _04720_ _02580_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_101_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_145_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput190 net190 la_data_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_98_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10073_ _04667_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09017__I _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06750__A1 net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10975_ _05407_ _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06502__A1 _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09687__I _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__I _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07058__A2 _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08255__B2 net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09598__A4 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11527_ _00311_ clknet_leaf_72_wb_clk_i net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_87_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _00242_ clknet_leaf_42_wb_clk_i as2650.PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_91_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10409_ _04882_ _04978_ _04980_ _04981_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_61_1827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_91_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11389_ _00015_ clknet_leaf_65_wb_clk_i as2650.cycle\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i clknet_4_12__leaf_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09507__A1 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05950_ _00943_ _00947_ _00950_ _00954_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__10117__A2 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05881_ _00887_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05919__I1 _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07620_ wb_counter\[20\] _02404_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07551_ _02341_ _02350_ _02352_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_85_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11192__I _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06502_ _01257_ _01460_ _01463_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_88_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06286__I _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07482_ _02237_ _02301_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09221_ _03886_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06433_ _01367_ _01395_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_4_13__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09038__A3 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09152_ _03679_ _03675_ _03645_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_115_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06364_ _01320_ _01328_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_40_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08103_ _02801_ _01892_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08797__A2 _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09083_ _03772_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06295_ _01266_ _01190_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_163_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08034_ _02788_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput70 net384 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput81 net412 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_9_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput92 net417 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08549__A2 _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__I _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09985_ _01835_ _04603_ _04606_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10271__I _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08936_ _01491_ _03584_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_122_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10108__A2 _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08867_ _03099_ _03559_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07818_ _02586_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07580__I _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08798_ as2650.stack\[12\]\[9\] _02533_ _02536_ as2650.stack\[13\]\[9\] _03494_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_168_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_8_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07749_ _02517_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output115_I net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06196__I _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _05214_ _05222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10292__A1 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09419_ _04094_ _04104_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_3_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10691_ _05168_ _05180_ _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_33_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08344__C _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11312_ _00108_ clknet_leaf_102_wb_clk_i net279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_147_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11243_ _00039_ clknet_leaf_40_wb_clk_i as2650.stack\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10347__A2 _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07212__A2 _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11174_ as2650.stack\[13\]\[14\] _05542_ _05545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10125_ _04701_ _04703_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10056_ _01939_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_166_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_100_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08476__A1 _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10958_ _05290_ _00725_ _01525_ _05010_ _05291_ _05393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__09673__B1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_80_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10283__A1 _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_80_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10889_ _04314_ _04315_ _05312_ _05329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_156_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08228__A1 _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06834__I as2650.debug_psl\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08228__B2 net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10586__A2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06080_ net249 _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
Xhold106 wbs_dat_i[15] net452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold117 wbs_dat_i[16] net463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_106_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_78_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08400__A1 _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08951__A2 _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09770_ _04450_ _04452_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06982_ _01742_ _01893_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_33_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05765__A2 _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06962__A1 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08721_ _01846_ _03351_ _03416_ _03059_ _03419_ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05933_ _00784_ _00810_ _00934_ _00937_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_87_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09900__A1 _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ as2650.stack\[0\]\[4\] _03302_ _03303_ as2650.stack\[1\]\[4\] _03294_ _03353_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05864_ _00689_ _00870_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07603_ net381 _02394_ _02385_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _00606_ _00610_ _03269_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05795_ _00804_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_136_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07534_ _02321_ _02337_ _02338_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08467__A1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10274__A1 _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07465_ _02278_ wb_counter\[28\] _02272_ _02287_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09204_ _03886_ _03887_ _03889_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_92_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08219__A1 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06416_ _01343_ _01379_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_27_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06744__I _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07396_ net274 _02225_ _02218_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09135_ _01281_ _01166_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06347_ as2650.cycle\[1\] _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_161_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09066_ _03754_ _03747_ _02482_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_128_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06278_ _01249_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_1834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06245__A3 _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08017_ _02771_ _02751_ _02772_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09719__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09968_ _04594_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08919_ _00828_ _01226_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09899_ _03153_ _02475_ _04551_ _04552_ as2650.trap _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__07524__B _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06919__I _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05823__I net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11861_ net299 net263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10812_ _05112_ _05249_ _05254_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11792_ _00571_ clknet_leaf_110_wb_clk_i as2650.stack\[13\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10743_ as2650.stack\[8\]\[14\] _05209_ _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10674_ _05171_ _05167_ _05170_ _00867_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_165_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10017__A1 as2650.stack\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09958__A1 _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05819__I0 _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06236__A3 _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11226_ _00022_ clknet_leaf_17_wb_clk_i as2650.stack\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08933__A2 _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11157_ _05457_ _05529_ _05534_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_156_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06944__A1 _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10740__A2 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10108_ as2650.stack\[3\]\[13\] _04688_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11088_ as2650.regs\[7\]\[6\] _05491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10039_ _01868_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_121_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06829__I _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_82_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_125_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_82_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05580_ _00593_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09646__B1 _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09110__A2 _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06564__I as2650.io_bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07250_ _02097_ _02083_ _02098_ _02099_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_119_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06201_ net54 _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09949__A1 as2650.io_bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07181_ _02045_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10559__A2 _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06132_ _00671_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold106_I wbs_dat_i[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06063_ as2650.PC\[0\] _00641_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05825__I3 _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05908__I _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09177__A2 _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _04329_ _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08924__A2 _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06935__A1 _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09753_ _01874_ _01102_ _04436_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06965_ _01877_ _01862_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XANTENNA__09543__C _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08704_ _01574_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05916_ _00753_ _00920_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09684_ _02562_ _04369_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_158_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06896_ _01812_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__05643__I as2650.cycle\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08635_ _01443_ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05847_ _00854_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_167_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08566_ _00606_ _03269_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05778_ _00689_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_77_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10247__A1 _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07517_ _02091_ wb_counter\[1\] _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05799__B _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ as2650.stack\[0\]\[0\] _02525_ _02528_ as2650.stack\[1\]\[0\] _02504_ _03202_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_65_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06474__I _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07448_ _02082_ wb_counter\[25\] _02270_ _02273_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_0_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A1 _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07379_ _02183_ _01560_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09118_ _03701_ _03705_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07415__A2 _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output182_I net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _04963_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_81_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09049_ _01411_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05977__A2 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10970__A2 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11011_ _01694_ _05186_ _04665_ _05437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_165_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08915__A2 _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06926__A1 _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_161_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09340__A2 _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10238__A1 _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11775_ _00554_ clknet_leaf_116_wb_clk_i as2650.stack\[14\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__A3 _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold84_I wbs_we_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06384__I _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10726_ _05092_ _05196_ _05201_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08851__B2 as2650.stack\[13\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10657_ _04931_ _05156_ _05157_ _04938_ _05158_ _05159_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_TAPCELL_ROW_114_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06209__A3 _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10588_ _01958_ _05112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_51_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10410__A1 _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10634__I _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08906__A2 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11209_ as2650.stack\[9\]\[11\] _05563_ _05567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07943__I _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10713__A2 _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06393__A2 _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ net252 _01617_ _01600_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_69_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05701_ _00680_ _00698_ _00713_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06681_ _01603_ _01609_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06145__A2 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07342__A1 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08420_ as2650.stack\[12\]\[15\] _02534_ _02537_ as2650.stack\[13\]\[15\] _03140_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05632_ _00645_ as2650.extend _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10229__A1 _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ _02765_ _03072_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09095__A1 _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07302_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06294__I as2650.relative_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08282_ _03000_ _02608_ net205 _03002_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_15_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05656__A1 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_60_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07233_ _02064_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_73_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_93_wb_clk_i clknet_4_10__leaf_wb_clk_i clknet_leaf_93_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_14_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07164_ _02035_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_22_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_22_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_30_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06115_ _01087_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_28_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07095_ as2650.stack\[11\]\[10\] _01987_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08070__A2 _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05638__I as2650.instruction_args_latch\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06081__A1 net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08014__I _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06046_ _01030_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_58_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06908__A1 _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_54_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input39_I io_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ _02557_ _04485_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07997_ _02627_ _02644_ _02753_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09736_ _01565_ _03714_ _04420_ _02562_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06948_ _01861_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_2_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09667_ _03768_ _04352_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06879_ _01795_ _01706_ _01796_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11649__CLK clknet_4_10__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06136__A2 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ _03317_ _03320_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07884__A2 _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09598_ _01674_ _01418_ _01648_ _01615_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_16_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05895__A1 net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08549_ as2650.stack\[0\]\[1\] _03249_ _03251_ as2650.stack\[1\]\[1\] _03252_ _03253_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_49_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11560_ _00344_ clknet_leaf_89_wb_clk_i as2650.stack\[10\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10511_ _04643_ _05053_ _05058_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11491_ _00275_ clknet_leaf_15_wb_clk_i as2650.stack\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_150_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10442_ _04156_ _04782_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05662__A4 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10373_ _03856_ _04808_ _04744_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07249__B _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_163_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09010__A1 _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06379__I _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_103_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_64_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11758_ _00537_ clknet_leaf_97_wb_clk_i as2650.regs\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_116_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10709_ as2650.stack\[8\]\[0\] _05191_ _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11689_ _00473_ clknet_leaf_114_wb_clk_i as2650.stack\[8\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11187__A2 _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ _02679_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09001__A1 _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08769__I _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09552__A2 _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ _02616_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_140_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_140_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_1656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06802_ as2650.is_interrupt_cycle _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 bus_in_gpios[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07782_ _02550_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09521_ _03689_ _03841_ _04206_ _02920_ _03842_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_79_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06733_ _01656_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09304__A2 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09452_ _04136_ _04137_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06664_ _01593_ _01591_ _01595_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08403_ _03036_ _03099_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05615_ as2650.indirect_target\[11\] _00626_ _00628_ as2650.PC\[11\] _00629_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_4_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09383_ net354 _04067_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10870__A1 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09068__A1 _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06595_ _01542_ net176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08334_ _02723_ _03055_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08009__I _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08265_ as2650.instruction_args_latch\[7\] _02975_ _02995_ _02981_ _02996_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08291__A2 _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__I _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07216_ _02070_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06752__I _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _01261_ _01298_ _01324_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_63_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_127_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ _02026_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_89_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09240__A1 _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07784__S _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10207__C _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07078_ _01801_ _01973_ _01979_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06029_ _01018_ net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_80_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10689__A1 _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_98_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09719_ _02590_ _02567_ _02991_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10991_ _02201_ as2650.regs\[4\]\[4\] _02669_ _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__07157__I1 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07306__A1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11102__A2 _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06927__I _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09059__A1 _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11612_ _00396_ clknet_leaf_130_wb_clk_i as2650.stack\[1\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06380__I2 net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10613__A1 _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11543_ _00327_ clknet_leaf_117_wb_clk_i as2650.stack\[4\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__A2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__I _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11474_ _00258_ clknet_leaf_30_wb_clk_i as2650.debug_psu\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10184__I _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10425_ _04849_ _04993_ _04996_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_1458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10356_ _04929_ _04930_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_143_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07793__A1 _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i clknet_4_11__leaf_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10287_ _04754_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06060__A4 _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__A2 _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A2 _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09298__B2 _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07148__I1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05741__I as2650.debug_psl\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06520__A2 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06380_ _00787_ net192 net201 _01025_ _01186_ _01188_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_139_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08273__A2 _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08050_ _02794_ _02799_ _02804_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06572__I _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10308__B _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07001_ _01904_ _01911_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_109_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10094__I _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10907__A2 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06426__I3 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08952_ _03619_ _03621_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08499__I _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07903_ _01170_ _01300_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08883_ _01934_ _03283_ _03241_ _03575_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_100_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06339__A2 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07834_ _02601_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_1586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_95_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07765_ _02533_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09551__C _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07139__I1 net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09828__A3 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06716_ _01640_ _01348_ _01641_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09504_ _03736_ _03416_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07839__A2 _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07696_ _01577_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09435_ _04093_ _04105_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10843__A1 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06647_ as2650.chirp_ptr\[0\] _01580_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_47_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09366_ _01029_ _01017_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06578_ _01077_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_1_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08317_ _03021_ _02803_ _03022_ net211 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_117_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09297_ _00825_ _00888_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_118_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08248_ as2650.instruction_args_latch\[4\] _02975_ _02980_ _02981_ _02982_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08179_ _01292_ _01305_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08016__A2 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10210_ _04724_ _04768_ _04771_ _04785_ _04787_ _04788_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_31_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11190_ _05447_ _05549_ _05555_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08567__A3 _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10141_ _01728_ _04717_ _04718_ _04719_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_24_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput180 net180 io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput191 net191 la_data_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10072_ _04666_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_140_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10126__A3 _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09742__B _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10974_ _02201_ _05286_ _05407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_134_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09033__I _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10179__I _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__A2 _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08255__A2 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10062__A2 _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11526_ _00310_ clknet_leaf_73_wb_clk_i net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_41_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_134_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11457_ _00241_ clknet_leaf_36_wb_clk_i as2650.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_145_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10408_ _01423_ _04758_ _04898_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_91_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11388_ _00014_ clknet_leaf_66_wb_clk_i as2650.cycle\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06569__A2 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10339_ _01656_ _04808_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07437__B _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07518__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10117__A3 _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08715__B1 _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05880_ as2650.regs\[1\]\[2\] as2650.regs\[5\]\[2\] _00800_ _00887_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07550_ net101 _02344_ _02351_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06501_ _01183_ _01461_ _01462_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_92_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07481_ net290 _02238_ _02300_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09691__A1 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08494__A2 _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09878__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09220_ _03904_ _03905_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_75_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06432_ _01347_ _01376_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_130_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09151_ _03675_ _03645_ _03679_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08715__C _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06363_ _01261_ _01327_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08102_ _02787_ _01907_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09082_ _01698_ _01280_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_66_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06294_ as2650.relative_cyc _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_86_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08033_ _02787_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput60 rom_bus_in[2] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_128_1475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput71 net426 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput82 net413 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput93 net391 net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_38_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09984_ as2650.stack\[4\]\[5\] _04604_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_1637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _03625_ _03626_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_157_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08866_ _03030_ _03098_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08182__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input21_I bus_in_sid[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07861__I _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07817_ _02585_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08797_ as2650.stack\[8\]\[9\] _02492_ _02499_ as2650.stack\[9\]\[9\] _02505_ _03493_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_93_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07748_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07679_ net248 net238 _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output108_I net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06496__A1 _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09418_ _04098_ _04103_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_133_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10690_ _05180_ _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10727__I _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09349_ _04033_ _04034_ _04026_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__06248__A1 _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11311_ _00107_ clknet_leaf_105_wb_clk_i net278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11242_ _00038_ clknet_leaf_15_wb_clk_i as2650.stack\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07257__B _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11173_ _05473_ _05541_ _05544_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06420__A1 _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10124_ _04702_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10055_ _04653_ _04646_ _04654_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07771__I _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08173__A1 _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_123_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06387__I net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09673__A1 _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08476__A2 _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10957_ as2650.regs\[4\]\[7\] _05335_ _05392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09673__B2 _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10888_ _05320_ _05327_ _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_1739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08228__A2 _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__A1 _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__A2 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11509_ _00293_ clknet_leaf_69_wb_clk_i net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_83_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold107 wbs_dat_i[20] net453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_41_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold118 wbs_dat_i[1] net464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_106_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06850__I _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08400__A2 _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06411__A1 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06981_ _01892_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_33_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05932_ _00770_ _00936_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_33_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08720_ _03284_ _03418_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_47_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08164__A1 _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08651_ as2650.stack\[3\]\[4\] _03289_ _03296_ as2650.stack\[2\]\[4\] _03352_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05863_ as2650.regs\[0\]\[1\] _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07911__A1 as2650.wb_hidden_rom_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07602_ _02339_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_59_1598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08582_ _01789_ _03270_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05794_ _00788_ _00794_ _00799_ _00803_ _00735_ _00768_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_77_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07533_ net358 _02323_ _02330_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09664__A1 as2650.debug_psl\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08726__B _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06478__A1 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07464_ net109 _02279_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_147_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06415_ _01344_ _01378_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_27_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09203_ _03888_ _00914_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07395_ _02211_ wb_counter\[17\] _02228_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09134_ _03752_ _03821_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06346_ _01312_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09065_ _03755_ _03268_ _03723_ net199 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06277_ as2650.cycle\[4\] _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_32_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08016_ _02625_ _01815_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ _01694_ _01713_ _04523_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06953__A2 _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08918_ _03607_ _03609_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_99_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07591__I _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09898_ _02559_ _03403_ _01228_ _04551_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA_output225_I net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08849_ as2650.stack\[11\]\[11\] _03141_ _01968_ as2650.stack\[10\]\[11\] _03543_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11860_ net171 net262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_1832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10811_ as2650.stack\[6\]\[15\] _05250_ _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11791_ _00570_ clknet_leaf_110_wb_clk_i as2650.stack\[13\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09655__A1 _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10742_ _05108_ _05208_ _05211_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10673_ _04834_ _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_54_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_24_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07969__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05819__I1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08630__A2 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06641__A1 _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06670__I _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11225_ _00021_ clknet_leaf_16_wb_clk_i as2650.stack\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09981__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11156_ as2650.stack\[13\]\[7\] _05530_ _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _04655_ _04687_ _04689_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_125_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11087_ _05177_ _05487_ _05488_ _05490_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_125_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10038_ _04641_ _04636_ _04642_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_121_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06200_ as2650.insin\[4\] _01096_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11205__A1 as2650.stack\[9\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10008__A2 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07180_ net87 net119 _02041_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06131_ _00669_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06062_ _01043_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06580__I _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08385__A1 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09821_ _04500_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10830__I _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ net188 _02473_ _04435_ _01275_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06964_ as2650.PC\[8\] _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08703_ _03344_ _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_154_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05915_ as2650.regs\[0\]\[4\] _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09683_ _04293_ _04302_ _04304_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06895_ as2650.PC\[4\] _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05846_ _00853_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_08634_ _00602_ _03285_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_90_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05777_ _00787_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09637__A1 as2650.debug_psu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ _01720_ _01128_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10247__A2 _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07516_ wb_counter\[0\] _02321_ _02324_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09101__A3 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08496_ as2650.stack\[3\]\[0\] _03200_ _02511_ as2650.stack\[2\]\[0\] _03201_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_130_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07447_ _02271_ _02272_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_130_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08860__A2 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05674__A2 _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07378_ net128 _02199_ _02213_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06329_ _01297_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09117_ _03753_ _03805_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08612__A2 _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11578__CLK clknet_leaf_92_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06490__I _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06623__A1 as2650.insin\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ _03698_ _03725_ _03734_ _03739_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_103_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output175_I net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10970__A3 _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11010_ _01736_ _05436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_165_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10183__A1 _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_161_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08128__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_1440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10486__A2 _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09628__A1 _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11774_ _00553_ clknet_leaf_111_wb_clk_i as2650.stack\[14\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07103__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09041__I _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10725_ as2650.stack\[8\]\[7\] _05197_ _05201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08851__A2 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_109_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10656_ as2650.regs\[1\]\[4\] _05159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_114_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_114_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10587_ _05110_ _05105_ _05111_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09800__A1 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_75_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06090__A2 net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08367__A1 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11208_ _05465_ _05562_ _05566_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_118_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11139_ _05523_ _05524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05700_ _00706_ net203 _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_69_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06680_ _01604_ _01608_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__A2 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05631_ as2650.indirect_cyc _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08350_ net208 _01437_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06575__I _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07301_ _02009_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_127_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08281_ _01258_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_24_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07232_ _02056_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_55_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05656__A2 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07163_ _02013_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10825__I _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06114_ _01086_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_112_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07094_ _01899_ _01986_ _01989_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06045_ _01029_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_62_wb_clk_i clknet_4_12__leaf_wb_clk_i clknet_leaf_62_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_105_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08358__A1 _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10560__I _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _01701_ _04477_ _04484_ _04480_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_157_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05654__I net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _02647_ _02752_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09735_ _03709_ _01201_ _03717_ _04406_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06947_ _01844_ _01860_ _01827_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_138_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09666_ _04333_ _04349_ _04351_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08965__I _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06878_ _01708_ _01710_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08530__A1 _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08617_ _03128_ _03319_ _01548_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05829_ _00835_ _00837_ _00657_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09597_ _01637_ _01625_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08186__B _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05895__A2 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08548_ _02503_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_166_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_13_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07097__A1 as2650.stack\[11\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08479_ as2650.ivectors_base\[11\] _03180_ _03182_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10510_ as2650.stack\[1\]\[7\] _05054_ _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output292_I net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11490_ _00274_ clknet_leaf_2_wb_clk_i as2650.stack\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10441_ _01857_ _04932_ _05012_ _04876_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_150_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10372_ _04794_ _04943_ _04945_ _04731_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_167_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i clknet_4_10__leaf_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_163_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08349__A1 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10470__I _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05583__A1 _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_1444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11757_ _00536_ clknet_leaf_97_wb_clk_i as2650.regs\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_116_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08824__A2 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10708_ _05190_ _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10631__A2 _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11688_ _00472_ clknet_leaf_114_wb_clk_i as2650.stack\[8\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10639_ _05145_ _05146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_153_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06063__A2 _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07260__A1 _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07012__A1 _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ _02615_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_120_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06801_ _00645_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07781_ _02549_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput3 bus_in_gpios[2] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09520_ _01703_ _04205_ _03688_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06732_ _00805_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06118__A3 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09451_ net218 net193 _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06663_ _01593_ _01587_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_135_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05614_ _00623_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08402_ _03036_ _02905_ _03099_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06594_ _01538_ _01514_ _01541_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_0_34_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09382_ _04067_ _04059_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_148_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_163_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08333_ _02934_ _03054_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08815__A2 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08264_ _01259_ _02993_ _02994_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06826__A1 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07215_ net159 net72 _02069_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08195_ _01265_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08579__A1 _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07146_ net102 net136 _02025_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08025__I _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10386__A1 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_144_Left_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07077_ as2650.stack\[11\]\[3\] _01975_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I ram_bus_in[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07864__I _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06028_ _01017_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_1657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output138_I net138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07979_ as2650.indirect_target\[3\] _02724_ _02735_ _02736_ _02737_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_138_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09718_ _03799_ _04402_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10990_ _05408_ _05419_ _05420_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07306__A2 _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_153_Left_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09649_ _02827_ _01669_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10310__B2 _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_156_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11611_ _00395_ clknet_leaf_129_wb_clk_i as2650.stack\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06380__I3 _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11542_ _00326_ clknet_leaf_126_wb_clk_i as2650.stack\[4\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06943__I _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_1436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11473_ _00257_ clknet_leaf_30_wb_clk_i as2650.debug_psu\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_162_Left_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10424_ _04853_ _04995_ _04731_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10377__A1 _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07242__A1 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10355_ _03847_ _04844_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10286_ _04860_ _04862_ _04756_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_109_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_105_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_66_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09298__A2 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07215__S _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10301__A1 _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_17_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_1549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10852__A2 _05282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07014__I _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06520__A3 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07949__I _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06853__I _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07481__A1 net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10375__I _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07000_ _01849_ _01909_ _01910_ _01842_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_96_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08951_ _03640_ _03642_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_102_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_51_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07902_ _02632_ _02652_ _02663_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08882_ _01936_ _03375_ _03574_ _03242_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08733__B2 as2650.stack\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ _00681_ _00685_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_93_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ _02532_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09503_ _04187_ _04188_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_155_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06715_ _01605_ _01501_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07695_ _01101_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_49_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09434_ _04117_ _04119_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06646_ _01582_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10843__A2 _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09365_ _04015_ _04049_ _04050_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06577_ _01525_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08464__B _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07859__I _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08316_ _03039_ _03040_ _03028_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09296_ _00766_ _01019_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _01001_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07472__A1 net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08178_ _02895_ _02917_ _02922_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_127_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07129_ _02016_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11020__A2 _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10140_ _01695_ _02917_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_28_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output255_I net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 net170 io_oeb[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput181 net306 io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput192 net192 la_data_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10071_ _01961_ _01970_ _04665_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08724__A1 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06938__I _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10973_ _05282_ _05398_ _05402_ _05406_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_85_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06502__A3 _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11525_ _00309_ clknet_leaf_72_wb_clk_i net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_134_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11456_ _00240_ clknet_leaf_43_wb_clk_i as2650.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10407_ _03857_ _04818_ _04979_ _04814_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_111_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11387_ _00013_ clknet_leaf_54_wb_clk_i as2650.cycle\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_91_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08963__A1 _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10338_ _04795_ _04911_ _04912_ _04801_ _00923_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_10__leaf_wb_clk_i clknet_leaf_119_wb_clk_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10269_ _04845_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_128_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05919__I3 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_85_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06500_ _01283_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07480_ _02094_ _02298_ _02299_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_92_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09691__A2 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06431_ _01393_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_44_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05701__A1 _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_98_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06362_ _01321_ _01322_ _01326_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09150_ _03823_ _03680_ _03836_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_98_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10589__A1 as2650.stack\[15\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08101_ _01002_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_40_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06293_ _01264_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08651__B1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09081_ _03694_ _03654_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08032_ _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_71_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput50 ram_bus_in[0] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput61 rom_bus_in[3] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput72 net420 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09827__C _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput83 net418 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_102_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput94 net416 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__A1 _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08303__I _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05768__A1 _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09983_ _01820_ _04603_ _04605_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08934_ _01497_ _01620_ _03584_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08706__B2 as2650.stack\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08865_ _02674_ _03555_ _03558_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_140_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07816_ _01233_ _01513_ _02583_ _02584_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_165_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_169_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08796_ as2650.stack\[11\]\[9\] _02509_ _02512_ as2650.stack\[10\]\[9\] _03492_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input14_I bus_in_serial_ports[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07747_ as2650.debug_psu\[2\] _02515_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_95_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_154_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09131__A1 _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10816__A2 _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07678_ _01055_ _01552_ _02451_ _02453_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_36_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09417_ _04099_ _04102_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06629_ _01556_ _01567_ _01571_ net179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09348_ _01495_ _01018_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ _03963_ _03964_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11310_ _00106_ clknet_leaf_140_wb_clk_i net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_50_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11241_ _00037_ clknet_leaf_15_wb_clk_i as2650.stack\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05759__A1 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ as2650.stack\[13\]\[13\] _05542_ _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_1705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10123_ _02714_ _01279_ _01508_ _02581_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_10054_ as2650.stack\[10\]\[11\] _04647_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10504__A1 as2650.stack\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08173__A2 _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05931__A1 _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_1633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10807__A2 _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10956_ _04313_ _05263_ _05390_ _05391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__09673__A2 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07684__A1 net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08881__B1 _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10887_ _04231_ _05276_ _05325_ _05326_ _05327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_136_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09425__A2 _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11508_ _00292_ clknet_leaf_67_wb_clk_i net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_129_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold108 wbs_dat_i[25] net454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__10991__A1 _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold119 wbs_dat_i[23] net465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_11439_ _00223_ clknet_leaf_60_wb_clk_i as2650.insin\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08936__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_1384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06980_ _01890_ _01891_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input6_I bus_in_gpios[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05931_ _00744_ as2650.instruction_args_latch\[7\] _00749_ _00935_ _00936_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_33_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08279__B _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08650_ _03288_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05862_ _00869_ net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10321__C _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07601_ wb_counter\[17\] _02392_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_55_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07911__A2 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ _01444_ _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_87_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_87_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05793_ _00800_ as2650.regs\[4\]\[5\] _00802_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_156_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07532_ _02131_ _02336_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_7_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_16_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_16_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07463_ _02277_ _02285_ _02286_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08872__B1 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09202_ _01023_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06414_ _01346_ _01377_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07394_ _02192_ _01874_ _02227_ _02170_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_17_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ _03753_ _03815_ _03820_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06345_ as2650.cycle\[2\] _01290_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08624__B1 _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06276_ _01241_ _01247_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09064_ _03754_ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05989__A1 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10982__A1 _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08015_ _02625_ _01815_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10563__I _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05657__I _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08033__I _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09966_ _01488_ _01675_ _04593_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08917_ _00923_ _03586_ _03608_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09897_ _03158_ _01285_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08848_ _03538_ _03539_ _03540_ _03541_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_output120_I net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output218_I net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08779_ _03337_ _03460_ _03475_ _03058_ _01307_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09104__A1 _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10810_ _05110_ _05249_ _05253_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11790_ _00569_ clknet_leaf_110_wb_clk_i as2650.stack\[13\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09655__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07666__A1 net400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10738__I _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10741_ as2650.stack\[8\]\[13\] _05209_ _05211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10672_ _05163_ _05167_ _05170_ _00848_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_24_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11214__A2 _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05819__I2 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A1 _05282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10406__C _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11224_ _00020_ clknet_leaf_2_wb_clk_i as2650.stack\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_112_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09591__A1 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11155_ _05455_ _05529_ _05533_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07782__I _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold22_I net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10106_ as2650.stack\[3\]\[12\] _04688_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_125_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11086_ as2650.regs\[7\]\[5\] _05490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_95_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10422__B _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10037_ as2650.stack\[10\]\[6\] _04637_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10141__C _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05904__A1 _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07657__A1 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10939_ _05315_ _04984_ _05374_ _05375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_27_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07022__I as2650.debug_psu\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09658__B _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08606__B1 _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06130_ as2650.extend _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06861__I as2650.debug_psl\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08082__A1 _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_134_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_134_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06061_ _00859_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_124_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__A1 _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09820_ _03105_ _04499_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08385__A2 _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06396__A1 _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09751_ _02484_ _04434_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06963_ _01874_ _01731_ _01875_ _01840_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_146_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08702_ _03343_ _01846_ _03240_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_94_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05914_ net200 _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06148__A1 _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09682_ _02583_ _03699_ _03799_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07196__I0 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06894_ _01804_ _01805_ _01810_ _01783_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08633_ _03329_ _03334_ _03267_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_90_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05845_ _00715_ as2650.regs\[4\]\[0\] _00852_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_08564_ _03258_ _03266_ _03267_ _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_49_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05776_ _00693_ _00785_ _00786_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_76_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07648__A1 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07515_ net72 _02323_ _02293_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08845__B1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08495_ _01689_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_159_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07446_ _02067_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_21_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07377_ _02121_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08472__B _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09116_ _03403_ _03803_ _03804_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06328_ _01296_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08073__A1 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06771__I _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10955__A1 _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06623__A2 wb_debug_cc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09047_ _03706_ _03737_ _03725_ _03738_ _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07820__A1 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06259_ _01206_ _01229_ _01231_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_108_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09573__A1 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09949_ as2650.io_bus_we _04554_ _04584_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_161_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08128__A2 _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09325__A1 _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06139__A1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07187__I0 net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05898__B1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09089__B1 _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11773_ _00552_ clknet_leaf_116_wb_clk_i as2650.stack\[14\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08300__A2 as2650.instruction_args_latch\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10724_ _05090_ _05196_ _05200_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10655_ _05150_ _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_84_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08064__A1 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ as2650.stack\[15\]\[14\] _05106_ _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_114_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10946__A1 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09800__A2 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11207_ as2650.stack\[9\]\[10\] _05563_ _05566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09564__A1 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10174__A2 as2650.instruction_args_latch\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11138_ _05520_ _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_78_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_4_15__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11069_ _00180_ _01594_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07178__I0 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11123__A1 as2650.stack\[14\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05630_ as2650.page_reg\[2\] _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_118_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07300_ _02130_ _02144_ _02145_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_24_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _02846_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07231_ _02081_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_6_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08292__B _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold111_I wbs_dat_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07162_ _02034_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06113_ _01085_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07093_ as2650.stack\[11\]\[9\] _01987_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06044_ _01028_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08358__A2 _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06369__A1 _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09803_ _02475_ _04483_ _02665_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08311__I _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07030__A2 _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07995_ _02626_ _01815_ _02751_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__09307__A1 _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _04291_ _04313_ _04418_ _02944_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06946_ as2650.PC\[7\] _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07169__I0 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11114__A1 _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_wb_clk_i clknet_4_6__leaf_wb_clk_i clknet_leaf_31_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_2_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07869__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09665_ _01754_ _04333_ _04350_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_2_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06877_ _01238_ _01243_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_59_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ _03082_ _03318_ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08530__A2 _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05828_ net305 _00836_ _00612_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09596_ _01383_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06392__I1 _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08547_ _03250_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05759_ _00748_ as2650.instruction_args_latch\[6\] _00749_ _00769_ _00770_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_132_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08478_ _00774_ _03179_ _03184_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07429_ net118 _02168_ _02150_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_4_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10440_ _03146_ _04934_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output285_I net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_167_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09794__A1 _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10371_ _04803_ _04944_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_167_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08349__A2 _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11756_ _00535_ clknet_leaf_94_wb_clk_i as2650.regs\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10707_ _05187_ _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11687_ _00471_ clknet_leaf_114_wb_clk_i as2650.stack\[8\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08037__A1 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10638_ _04695_ _05144_ _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_49_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10919__A1 _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10569_ as2650.stack\[15\]\[9\] _05096_ _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09537__A1 _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06800_ _01720_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07780_ _02548_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_1669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 bus_in_gpios[3] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06731_ _01648_ _01601_ _01655_ net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_116_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06118__A4 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09450_ _00721_ _00767_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06662_ _01593_ _01594_ _01590_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06523__A1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ _03106_ _03121_ _02667_ _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05613_ as2650.indirect_target\[10\] _00626_ _00623_ as2650.PC\[10\] _00627_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_56_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09381_ _04061_ _04063_ _04066_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_06593_ _01003_ _01306_ _01539_ _01540_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08332_ _02636_ _00958_ _03053_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10083__A1 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08263_ as2650.instruction_args_latch\[7\] _02978_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07214_ _02062_ _02068_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_61_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08028__A1 as2650.ivectors_base\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ _02935_ _01202_ _01222_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ _02014_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_42_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07076_ _01777_ _01973_ _01978_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09565__C _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09528__A1 _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10571__I _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06027_ _01016_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input44_I irqs[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07978_ _01468_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_96_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07880__I _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09717_ _03769_ _04400_ _04401_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06929_ as2650.PC\[6\] _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09648_ _02813_ _01677_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output200_I net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09579_ net217 _01418_ _04264_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_1618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11610_ _00394_ clknet_leaf_128_wb_clk_i as2650.stack\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11541_ _00325_ clknet_leaf_137_wb_clk_i as2650.stack\[4\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08019__A1 _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11472_ _00256_ clknet_4_12__leaf_wb_clk_i as2650.debug_psl\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__A1 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10423_ _00738_ _04994_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_21_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _04927_ _04928_ _04831_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _04231_ _04861_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10129__A2 _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_168_Right_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06753__A1 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_17_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08258__A1 as2650.instruction_args_latch\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11808_ _00587_ clknet_leaf_111_wb_clk_i as2650.stack\[9\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11739_ _00523_ clknet_leaf_131_wb_clk_i as2650.stack\[0\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09758__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07965__I _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__B1 _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06441__B1 _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06587__A4 _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ _01212_ _01643_ _03641_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_122_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06992__A1 _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ as2650.indirect_target\[0\] _02654_ _02657_ _02662_ _02463_ _02663_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08881_ _03337_ _03562_ _03573_ _03324_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09930__A1 _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07832_ _02599_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07763_ _02490_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09502_ _01510_ _03151_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06714_ _01044_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07694_ _02462_ _01534_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_49_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08497__B2 as2650.stack\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09433_ _04098_ _04103_ _04118_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06645_ as2650.chirp_ptr\[2\] _01581_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_78_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09364_ _03985_ _01013_ _03893_ _00856_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_75_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06576_ _01515_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_164_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08315_ _03034_ _02895_ _03026_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_69_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09997__A1 _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09295_ _03972_ _03980_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_75_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08246_ _02968_ _02977_ _02979_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08036__I _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08177_ _02918_ _02921_ _02664_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_31_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07875__I _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07128_ net72 net122 _02015_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07224__A2 wb_feedback_delay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07059_ _01963_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput160 net160 cs_port[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput171 net171 io_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_output150_I net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput182 net182 io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput193 net193 la_data_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10070_ _02545_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output248_I net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10531__A2 _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10972_ as2650.regs\[0\]\[0\] _05405_ _05406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07115__I _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10295__A1 _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11860__I net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05849__I0 _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11524_ _00308_ clknet_leaf_73_wb_clk_i net222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_134_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11455_ _00239_ clknet_leaf_35_wb_clk_i as2650.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_145_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwire298 net186 net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_111_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_hold52_I net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07785__I _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10406_ _03036_ _01421_ _01420_ _04820_ _04819_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_33_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11386_ _00012_ clknet_leaf_66_wb_clk_i as2650.cycle\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_130_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10337_ _01505_ _04799_ _01397_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10268_ _01084_ _04380_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_1731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08715__A2 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10199_ _04777_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_128_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08549__C _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_21_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08479__A1 as2650.ivectors_base\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ _01360_ _01392_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09691__A3 _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06864__I _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09979__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06361_ _01325_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08100_ _02624_ _02851_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_40_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10589__A2 _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09080_ _03694_ _03690_ _03691_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06292_ _01263_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08031_ net64 _02763_ _02785_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xinput40 io_in[7] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput51 ram_bus_in[1] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput62 rom_bus_in[4] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_130_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput73 net372 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08403__A1 _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput84 net414 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 net399 net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_40_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__A2 _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10210__B2 _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09982_ as2650.stack\[4\]\[4\] _04604_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11010__I _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05768__A2 _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06104__I _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08933_ _03623_ _03624_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08864_ _03280_ _03552_ _03557_ _02657_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_140_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_140_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07815_ _01424_ _01508_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_77_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08795_ _03487_ _03488_ _03489_ _03490_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07746_ as2650.debug_psu\[0\] as2650.debug_psu\[1\] _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_168_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05940__A2 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09131__A2 _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ net228 _02452_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08475__B _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09416_ _04100_ _04101_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06628_ _01556_ _01570_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08890__A1 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09347_ _01500_ _04027_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06559_ _01001_ _01507_ _01513_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_118_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _00729_ _01017_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output198_I net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08229_ as2650.instruction_args_latch\[2\] _02955_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11240_ _00036_ clknet_leaf_157_wb_clk_i as2650.stack\[11\]\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10201__A1 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08945__A2 _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11171_ _05469_ _05541_ _05543_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05759__A2 as2650.instruction_args_latch\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10122_ _01502_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_101_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11855__I net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10053_ _01927_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06184__A2 _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05931__A2 as2650.instruction_args_latch\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10955_ _04365_ _05302_ _05388_ _05389_ _05312_ _05390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__08385__B _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07684__A2 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10886_ _04175_ _04781_ _05303_ _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_80_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11507_ _00291_ clknet_leaf_66_wb_clk_i net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__10440__A1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold109 wbs_dat_i[13] net455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_65_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11438_ _00222_ clknet_leaf_60_wb_clk_i as2650.insin\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11369_ _00165_ clknet_leaf_68_wb_clk_i net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__10743__A2 _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05930_ _00697_ _00720_ net203 _00729_ _00735_ _00768_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_119_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05861_ _00845_ _00867_ _00868_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06175__A2 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07600_ _02391_ _02387_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_156_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08580_ _01101_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05792_ _00715_ _00801_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_18_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10259__A1 _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07531_ _02335_ _02327_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_76_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07124__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07462_ net285 _02282_ _02275_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09201_ _00765_ _01013_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06413_ _01347_ _01376_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07393_ net113 _02168_ _02193_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_56_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09132_ _02573_ _03819_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06344_ _01311_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09063_ _03737_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06275_ _01246_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08014_ _02769_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_108_1826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08388__B1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08927__A2 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_5__f_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09965_ net227 _01545_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05610__B2 as2650.PC\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08916_ _03588_ _01651_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06769__I _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09896_ _01959_ _04545_ _04550_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08847_ as2650.stack\[4\]\[11\] _03137_ _03138_ as2650.stack\[5\]\[11\] _03117_ _03541_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06166__A2 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08778_ _03469_ _03474_ _03267_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09104__A2 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ _02497_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output113_I net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_7_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10740_ _05104_ _05208_ _05210_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07666__A2 _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10671_ _05169_ _05170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08652__C _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08918__A2 _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11223_ _00019_ clknet_leaf_2_wb_clk_i as2650.stack\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11154_ as2650.stack\[13\]\[6\] _05530_ _05533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09591__A2 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_4_13__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _04669_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11085_ _05174_ _05487_ _05488_ _05489_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_159_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10036_ _01852_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08551__B1 _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09004__B _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ _04364_ _04843_ _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10661__A1 _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10661__B2 _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10869_ _05303_ _05309_ _05310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_89_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09658__C _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10664__I _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06060_ _01040_ _01041_ _00749_ _00857_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_124_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08909__A2 _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07973__I _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10716__A2 _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_103_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_103_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06589__I _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06962_ net219 _01732_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09750_ _01874_ _04433_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08701_ _03107_ _02799_ _03399_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05913_ _00918_ net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09681_ _03716_ _04366_ _02562_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06893_ _01808_ _01809_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07196__I1 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08632_ _03330_ _03331_ _03332_ _03333_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05844_ _00753_ _00851_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08563_ _02549_ _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05775_ _00693_ as2650.regs\[7\]\[5\] _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09098__A1 _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07514_ _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_9_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08494_ _03158_ _01217_ _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_65_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07445_ _02010_ _02064_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10652__A1 _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10652__B2 _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07376_ _02115_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_21_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10404__A1 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09115_ _03733_ _03757_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06327_ _01171_ _01181_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10574__I _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08073__A2 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09046_ _03737_ _03218_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06258_ _01230_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_108_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08979__I _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06189_ _01097_ _01160_ _01161_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_44_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07883__I _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09573__A2 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ _04554_ _01529_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_161_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_161_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output230_I net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07336__A1 _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09879_ as2650.stack\[5\]\[8\] _04540_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07187__I1 net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_149_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_120_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05898__B2 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10749__I _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09089__A1 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11772_ _00551_ clknet_leaf_131_wb_clk_i as2650.stack\[14\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08836__A1 _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10723_ as2650.stack\[8\]\[6\] _05197_ _05200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10643__A1 _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05779__S _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_118_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10654_ _05148_ _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_118_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08382__C _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ _01953_ _05110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11520__D _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_1_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_75_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11206_ _05463_ _05562_ _05565_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11137_ _05521_ _05522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11068_ _05477_ _05470_ _05478_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07327__A1 net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07178__I1 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10019_ _01759_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_69_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05889__A1 _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10882__A1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08827__B2 _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__I _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07230_ _02066_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07161_ net78 net128 _02030_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08055__A2 _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10937__A2 _05369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06112_ _01084_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_hold104_I wbs_dat_i[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07092_ _01883_ _01986_ _01988_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05813__A1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06043_ _01027_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08799__I _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09802_ _01509_ _04476_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07994_ _02749_ _02729_ _02750_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09307__A2 _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06945_ _01857_ _01805_ _01858_ _01840_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09733_ _01856_ _03722_ _04416_ _04417_ _04291_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07169__I1 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09664_ as2650.debug_psl\[1\] _04334_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_39_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06876_ _01788_ _01793_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05827_ _00609_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08615_ _03077_ _03080_ _03081_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09595_ _03728_ _04280_ _03730_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
Xclkbuf_leaf_71_wb_clk_i clknet_4_12__leaf_wb_clk_i clknet_leaf_71_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_132_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08546_ _02496_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05758_ net211 _00758_ net202 _00767_ _00735_ _00768_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_72_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08477_ as2650.ivectors_base\[10\] _03180_ _03182_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09491__A1 _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05689_ _00702_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_163_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__I _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07428_ _02251_ _02255_ _02257_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07359_ net269 _02197_ _02188_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_1722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09243__A1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06057__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_149_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output180_I net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10370_ _01557_ _04282_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_167_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_167_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05804__A1 _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09029_ _03720_ _02471_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_14_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_163_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10864__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10479__I _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08809__A1 _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08285__A2 _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11755_ _00534_ clknet_leaf_95_wb_clk_i as2650.regs\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_165_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_hold82_I wbs_cyc_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10706_ _05188_ _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_165_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11686_ _00470_ clknet_leaf_127_wb_clk_i as2650.stack\[8\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10428__B _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10637_ _04698_ _04721_ _05143_ _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_24_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10568_ _01898_ _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08840__C _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10499_ _04631_ _05046_ _05051_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09508__I _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06730_ _01551_ _01653_ _01654_ _01612_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xinput5 bus_in_gpios[4] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07472__B _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_1372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06661_ _01589_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10389__I _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05612_ _00621_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08400_ _03107_ _03108_ _03120_ _03061_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09380_ _04048_ _04064_ _04065_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06592_ as2650.cycle\[2\] as2650.cycle\[8\] _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XANTENNA__09848__I0 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08331_ _03052_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10607__A1 _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07698__I _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05720__B _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ _01251_ _02992_ _02976_ net203 _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_117_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ _02010_ _02064_ _02065_ _02067_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__08028__A2 _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08193_ _01336_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11013__I _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07144_ _02024_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__A2 _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07787__A1 _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07075_ as2650.stack\[11\]\[2\] _01975_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06026_ _00866_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_125_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05893__S0 net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_58_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input37_I io_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06211__A1 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07977_ _02000_ _02734_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09716_ _02587_ _04365_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06928_ _01842_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_74_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09647_ _02812_ _01677_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06859_ as2650.stack\[12\]\[2\] _01739_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07711__A1 _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ _04254_ _04262_ _04263_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_156_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08529_ _02673_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09464__A1 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11540_ _00324_ clknet_leaf_137_wb_clk_i as2650.stack\[4\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07475__B1 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11471_ _00255_ clknet_leaf_87_wb_clk_i as2650.debug_psl\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _03855_ _01383_ _03580_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09767__A2 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11858__I net298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10353_ _04386_ _04846_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_76_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10284_ _04810_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10129__A3 _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06202__A1 _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07950__B2 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10837__A1 _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07702__A1 _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08608__S _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11807_ _00586_ clknet_leaf_111_wb_clk_i as2650.stack\[9\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10065__A2 _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ _00522_ clknet_leaf_24_wb_clk_i as2650.stack\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__I _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11669_ _00453_ clknet_leaf_94_wb_clk_i as2650.regs\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_94_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08430__A2 _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07900_ _02659_ _02661_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09682__B _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08880_ _03567_ _03572_ _02551_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07981__I _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08194__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07831_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07941__A1 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07762_ as2650.stack\[8\]\[13\] _02527_ _02530_ as2650.stack\[9\]\[13\] _02506_ _02531_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_75_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09501_ _01575_ _01578_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06713_ net242 net237 _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07693_ _01723_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09694__A1 as2650.cycle\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_49_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09432_ net218 net191 _04104_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06644_ as2650.chirp_ptr\[1\] as2650.chirp_ptr\[0\] _01580_ _01581_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_133_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06575_ _01524_ net157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09363_ _00817_ _03893_ _03938_ _03985_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_118_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08314_ _03029_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_151_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09294_ _03973_ _03979_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_75_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07221__I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08245_ as2650.instruction_args_latch\[4\] _02978_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11005__A1 _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08176_ _01130_ _02919_ _01206_ _02920_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__09749__A2 _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07127_ _02014_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_15_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10582__I _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_149_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07058_ _01872_ _01886_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_100_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput150 net150 bus_data_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08709__B1 _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput161 net161 cs_port[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06009_ _01008_ net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput172 net299 io_out[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput183 net183 io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput194 net194 la_data_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09921__A2 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06735__A2 _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _05404_ _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_1540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11523_ _00307_ clknet_4_15__leaf_wb_clk_i net236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_53_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06970__I _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11454_ _00238_ clknet_4_6__leaf_wb_clk_i as2650.PC\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire299 net172 net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_130_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10405_ _04976_ _04977_ _04750_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11385_ _00011_ clknet_leaf_55_wb_clk_i as2650.cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_130_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_1512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06423__A1 _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10336_ _01389_ _04798_ _04799_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_46_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10267_ _04763_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08176__A1 _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09912__A2 _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _01729_ _04188_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06210__I _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_128_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_128_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09691__A4 _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06366__B _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06360_ _01181_ _01324_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07439__B1 as2650.debug_psu\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09979__A2 _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08100__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_40_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06291_ _01262_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_4_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08030_ _01153_ _01145_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_167_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06880__I _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 bus_in_timers[5] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 io_in[8] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput52 ram_bus_in[2] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput63 rom_bus_in[5] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput74 net376 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput85 net419 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput96 net405 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_123_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06414__A1 _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10210__A2 _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09981_ _04597_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08932_ _02606_ _03583_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_62_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08167__A1 _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ _03020_ _03097_ _03556_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_122_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_140_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07814_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08794_ as2650.stack\[4\]\[9\] _02533_ _02536_ as2650.stack\[5\]\[9\] _02520_ _03490_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07745_ as2650.stack\[7\]\[13\] _02510_ _02513_ as2650.stack\[6\]\[13\] _02514_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_139_1596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09667__A1 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07676_ _01550_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09415_ _00757_ _03888_ _01029_ _00719_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10577__I _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06627_ _01569_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_94_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08890__A2 _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06558_ _01512_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08047__I _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09346_ _04030_ _04031_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06489_ _01314_ _01253_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_111_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09277_ _03949_ _03961_ _03962_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_62_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08642__A2 _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ _01252_ _02617_ _02952_ net197 _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_146_1545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _01949_ _01298_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_147_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11201__I _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10245__C _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11170_ as2650.stack\[13\]\[12\] _05542_ _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _03812_ _04699_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _04651_ _04646_ _04652_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10268__A2 _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10954_ _04168_ _04782_ _05303_ _05389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_84_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08330__A1 _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10885_ as2650.chirpchar\[2\] _05271_ _05324_ _05272_ _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_38_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09830__A1 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11506_ _00290_ clknet_leaf_66_wb_clk_i net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_136_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_94_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10991__A3 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11437_ _00221_ clknet_4_6__leaf_wb_clk_i as2650.page_reg\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11368_ _00164_ clknet_leaf_69_wb_clk_i net230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06947__A2 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10319_ _02894_ _01402_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08149__A1 _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11299_ _00095_ clknet_leaf_143_wb_clk_i net296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09960__B _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05860_ _00723_ as2650.regs\[6\]\[1\] _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05758__I0 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09649__A1 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ as2650.regs\[0\]\[5\] _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_37_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07530_ wb_counter\[3\] _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06875__I _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07124__A2 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07461_ _02278_ wb_counter\[27\] _02273_ _02284_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_134_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08872__A2 _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06412_ _00828_ _01375_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09200_ _00728_ _00889_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07392_ _02220_ _02224_ _02226_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05930__I0 _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06343_ as2650.cycle\[7\] _01290_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_112_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09131_ _03817_ _02628_ _03807_ _03818_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08624__A2 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06635__A1 _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09062_ _03703_ _03718_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06274_ as2650.cycle\[11\] _01245_ _01093_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10431__A2 _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_96_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_96_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05989__A3 _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08013_ _01160_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10982__A3 _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11021__I _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_25_wb_clk_i clknet_4_6__leaf_wb_clk_i clknet_leaf_25_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06115__I _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09964_ _01665_ _04592_ _01088_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08915_ _03605_ _03606_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09895_ as2650.stack\[5\]\[15\] _04546_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_139_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ as2650.stack\[7\]\[11\] _01692_ _01968_ as2650.stack\[6\]\[11\] _03540_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08777_ _03470_ _03471_ _03472_ _03473_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_154_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05989_ net224 _00956_ _00964_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_0_71_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07728_ _02496_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08312__B2 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07659_ wb_counter\[28\] _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output106_I net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10670__A2 _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10670_ _05168_ _05166_ _05169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ _00898_ _00889_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_24_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10422__A2 _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08505__I _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__A1 _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06641__A4 _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11222_ _00018_ clknet_leaf_2_wb_clk_i as2650.stack\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_112_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10186__A1 _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07051__A1 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11153_ _05453_ _05529_ _05532_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10104_ _04667_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11084_ as2650.regs\[7\]\[4\] _05489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_120_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09879__A1 as2650.stack\[5\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10035_ _04639_ _04636_ _04640_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_86_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07106__A2 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10937_ _05261_ _05369_ _05370_ _05373_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09004__C _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11106__I _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10010__I _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10868_ _05306_ _05307_ _05308_ _05309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08606__A2 _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09803__A1 _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10799_ as2650.stack\[6\]\[10\] _05244_ _05247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10949__B1 _05384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10680__I _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08790__A1 _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ _01873_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_24_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08700_ _02802_ _02642_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05912_ _00692_ _00916_ _00917_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09680_ _04364_ _04216_ _04249_ _04365_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_55_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06892_ _01752_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_143_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_143_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_136_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08631_ as2650.stack\[15\]\[3\] _03308_ _03142_ as2650.stack\[14\]\[3\] _03298_ _03333_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_94_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05843_ as2650.regs\[0\]\[0\] _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08562_ _03259_ _03260_ _03263_ _03265_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05774_ as2650.regs\[3\]\[5\] _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09098__A2 _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _02319_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08493_ _01219_ _01444_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08845__A2 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06856__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07444_ net121 _02119_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_58_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07375_ _02113_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_146_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09114_ _03755_ _03335_ _03723_ net214 _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06326_ _01294_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06257_ _01142_ _01165_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07281__A1 net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ _03736_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05831__A2 _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06188_ as2650.insin\[5\] _01097_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__A1 _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08060__I _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08781__B2 _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09947_ _02814_ _04578_ _04583_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__05595__A1 as2650.cycle\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09878_ _04527_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07336__A2 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output223_I net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08829_ as2650.stack\[8\]\[10\] _03261_ _03262_ as2650.stack\[9\]\[10\] _03464_ _03524_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_169_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10891__A2 _05330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11771_ _00550_ clknet_leaf_131_wb_clk_i as2650.stack\[14\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08836__A2 _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10722_ _05088_ _05196_ _05199_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10653_ _05145_ _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_165_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10584_ _05108_ _05105_ _05109_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_114_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07272__A1 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_71_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11205_ as2650.stack\[9\]\[9\] _05563_ _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07024__A1 _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11136_ _05520_ _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_97_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05586__A1 as2650.indirect_target\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11067_ as2650.stack\[0\]\[15\] _05471_ _05478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10018_ _04621_ _04625_ _04628_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10331__A1 _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_1728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06838__A1 _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10675__I _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07160_ _02033_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08145__I as2650.instruction_args_latch\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10398__A1 _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06111_ _01083_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_54_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06066__A2 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07091_ as2650.stack\[11\]\[8\] _01987_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06042_ _00922_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_105_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07015__A1 net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10343__C _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08763__A1 _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ _03502_ _04443_ _04479_ _04481_ _04439_ _03808_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
X_07993_ _02725_ _01791_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09732_ _03857_ _03731_ _03721_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06944_ _01565_ _01809_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_105_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09663_ _04334_ _04335_ _04338_ _04348_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_2_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06875_ _01785_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08614_ _02762_ _03282_ _03316_ _03278_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05826_ as2650.indirect_target\[3\] _00621_ _00623_ as2650.PC\[3\] _00835_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__10873__A2 _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09594_ _04279_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08545_ _03248_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06392__I3 _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05757_ _00704_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ _00794_ _03179_ _03183_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05688_ _00700_ _00681_ _00685_ _00701_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_108_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A2 _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07427_ net279 _02256_ _02249_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10585__I _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_114_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05679__I _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_40_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_40_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07358_ _02136_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06309_ as2650.insin\[5\] _01097_ _01279_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__07254__A1 net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07289_ _02077_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07894__I _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09028_ _02578_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output173_I net173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06303__I _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_123_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_156_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_107_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_103_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__A2 _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11754_ _00533_ clknet_leaf_79_wb_clk_i as2650.regs\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _05187_ _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07493__A1 net366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11685_ _00469_ clknet_leaf_21_wb_clk_i as2650.stack\[8\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10636_ _01807_ _05142_ _05143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_102_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07245__A1 net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _05094_ _05095_ _05097_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10498_ as2650.stack\[1\]\[2\] _05048_ _05051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08745__B2 _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11119_ as2650.stack\[14\]\[9\] _05509_ _05511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 bus_in_gpios[5] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06660_ _01592_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_153_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05611_ _00620_ _00622_ _00624_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_8_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06591_ _01142_ _01272_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_52_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08330_ _02683_ _01474_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06883__I _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07484__A1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08261_ _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08681__B1 _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _02056_ _02066_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08192_ _01249_ _01297_ _01302_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_85_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07143_ net101 net135 _02020_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09776__A3 _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07787__A2 _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07074_ _01760_ _01973_ _01977_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06025_ _01015_ net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_61_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09784__I0 _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06211__A2 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ _01326_ _02730_ _02733_ _02705_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_143_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09715_ _04399_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_143_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11099__A2 _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06927_ _01797_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_74_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09161__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09646_ _04305_ _04328_ _04331_ _03717_ _03769_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06858_ _01776_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05809_ _00707_ as2650.regs\[6\]\[3\] _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_156_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09577_ _01026_ _01656_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_156_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06789_ _01704_ _01709_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_78_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08528_ _03194_ _03196_ _03232_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_52_1755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09464__A2 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07475__A1 _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ _03162_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_1510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output290_I net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11470_ _00254_ clknet_leaf_83_wb_clk_i as2650.debug_psl\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10421_ _04795_ _04991_ _04992_ _04801_ _01856_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_85_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11023__A2 _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08424__B1 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10352_ _04924_ _04925_ _04926_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08513__I _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10782__A1 _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_1738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10283_ _01616_ _04848_ _04857_ _04859_ _04746_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XPHY_EDGE_ROW_131_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08727__A1 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10129__A4 _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06033__I _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05961__A1 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05713__A1 _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11806_ _00585_ clknet_leaf_111_wb_clk_i as2650.stack\[9\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07466__A1 net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11737_ _00521_ clknet_leaf_24_wb_clk_i as2650.stack\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11668_ _00452_ clknet_leaf_80_wb_clk_i as2650.regs\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10619_ _05098_ _05129_ _05132_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11599_ _00383_ clknet_leaf_122_wb_clk_i as2650.stack\[2\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07769__A2 _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08423__I _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10174__B _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06441__A2 _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07039__I _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08194__A2 _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ _02597_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05782__I _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07761_ _02529_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05952__A1 _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09500_ _04185_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06712_ _01550_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07692_ _01038_ _02452_ _02451_ _02461_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_155_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09694__A2 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09431_ _04115_ _04116_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06643_ _01574_ _01579_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_49_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09362_ _03888_ _01019_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_75_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06574_ as2650.io_bus_we _01519_ _01521_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_47_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08313_ _02935_ _02937_ _03036_ _03010_ _03037_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_111_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09293_ _03978_ _03977_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_74_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11024__I _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08244_ _02954_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06680__A2 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ _02564_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09749__A3 _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07126_ _02013_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07057_ _01901_ _01924_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xoutput140 net140 bus_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput151 net151 bus_data_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08709__A1 _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06008_ _00961_ _00994_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput162 net162 io_oeb[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput173 net173 io_out[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_105_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput184 net184 io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput195 net195 la_data_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_122_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07959_ _02462_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output136_I net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05794__I1 _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10970_ _04769_ _01515_ _05259_ _05403_ _05404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09629_ _01771_ _04307_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07448__A1 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07448__B2 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11522_ _00306_ clknet_leaf_73_wb_clk_i net235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07999__A2 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05849__I2 net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08671__C _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11453_ _00237_ clknet_leaf_35_wb_clk_i as2650.PC\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08948__A1 _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _04210_ _04811_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_130_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11384_ _00010_ clknet_leaf_49_wb_clk_i as2650.is_interrupt_cycle vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_91_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_91_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10335_ _03847_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_91_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10266_ _04763_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_20_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _03475_ _04775_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08418__I _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06290_ as2650.cycle\[6\] _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 bus_in_sid[3] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10683__I _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput31 bus_in_timers[6] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput42 io_in[9] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05777__I _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput53 ram_bus_in[3] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput64 rom_bus_in[6] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput75 net387 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput86 net425 net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput97 net365 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09980_ _04595_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08931_ _00881_ _01225_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11652__CLK clknet_leaf_92_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ _03098_ _03347_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_129_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07813_ _01204_ _01163_ _02581_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_140_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08793_ as2650.stack\[7\]\[9\] _02509_ _02512_ as2650.stack\[6\]\[9\] _03489_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09116__A1 _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07744_ _02512_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07678__A1 _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _01241_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08875__B1 _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09414_ _00718_ _03892_ _03888_ _01028_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06626_ _01568_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08328__I _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09345_ _04020_ _04022_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06557_ _01508_ _01511_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09276_ _03950_ _03951_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06488_ _01315_ _01331_ _01448_ _01449_ _01450_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__10985__A1 _05330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08227_ _02949_ _02963_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10593__I _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05687__I _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08158_ _00652_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_31_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07109_ _01307_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08089_ _02802_ _02825_ _02840_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05759__A4 _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10120_ _03159_ _04698_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output253_I net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10051_ as2650.stack\[10\]\[10\] _04647_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11162__A1 as2650.stack\[13\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07407__I _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07905__A2 _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06311__I _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05916__A1 _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09658__A2 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05931__A4 _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10953_ net194 _04773_ _05387_ _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_86_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06341__A1 _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10884_ _05322_ _05323_ _05304_ _05324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11217__A2 _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07141__I0 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11505_ _00289_ clknet_leaf_67_wb_clk_i net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_136_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_93_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11436_ _00220_ clknet_leaf_55_wb_clk_i as2650.page_reg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11367_ _00163_ clknet_leaf_69_wb_clk_i net229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_145_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10318_ _04892_ _04893_ _04750_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_123_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11298_ _00094_ clknet_leaf_144_wb_clk_i net295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08149__A2 _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10249_ _04790_ _04791_ _04816_ _04824_ _04826_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__11153__A1 _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09897__A2 _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05790_ as2650.debug_psl\[4\] _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_89_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09649__A2 _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07460_ net108 _02279_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_18_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06411_ _01371_ _01374_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07391_ net273 _02225_ _02218_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_1524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07987__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05930__I1 _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09130_ _03709_ _02627_ _02568_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06342_ _01310_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07132__I0 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10967__A1 _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09061_ _02003_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_66_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06635__A2 _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06273_ _01098_ _01244_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_142_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08012_ _02746_ _02747_ _02760_ _02768_ _02745_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__10346__C _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08388__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09585__A1 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09585__B2 _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09963_ net226 _04586_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_13__leaf_wb_clk_i clknet_leaf_65_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_141_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08914_ _01178_ _03585_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _01954_ _04545_ _04549_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08845_ as2650.stack\[0\]\[11\] _03137_ _03138_ as2650.stack\[1\]\[11\] _03131_ _03539_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_139_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08776_ as2650.stack\[15\]\[8\] _03244_ _03254_ as2650.stack\[14\]\[8\] _03256_ _03473_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05988_ net235 _00988_ _00974_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__05970__I _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06571__A1 as2650.io_bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I bus_in_serial_ports[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10588__I _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07727_ _02495_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08312__A2 _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07658_ _02423_ _02437_ _02438_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06609_ web_behavior\[1\] _01553_ clknet_leaf_149_wb_clk_i _01554_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_36_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07589_ wb_counter\[15\] _02382_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07897__I _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ _00914_ _01489_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09259_ _00756_ _00791_ _01493_ _03938_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__07823__A1 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11212__I _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__A2 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11221_ _00017_ clknet_leaf_3_wb_clk_i as2650.stack\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09576__A1 _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08521__I _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11152_ as2650.stack\[13\]\[5\] _05530_ _05532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09328__A1 _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10103_ _04653_ _04681_ _04686_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_1549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11083_ _05481_ _05488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_125_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10034_ as2650.stack\[10\]\[5\] _04637_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06041__I _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07581__B _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08551__A2 _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06562__A1 _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06909__C _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10936_ _05371_ _05372_ _05260_ _05373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06314__A1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10110__A2 _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10867_ _04038_ _04176_ _04963_ _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08067__B2 as2650.indirect_target\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10798_ _05098_ _05243_ _05246_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10166__C _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09567__A1 _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11419_ _00203_ clknet_leaf_71_wb_clk_i as2650.instruction_args_latch\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06960_ _01872_ _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07047__I _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I bus_in_gpios[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05911_ _00847_ as2650.regs\[6\]\[4\] _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06891_ _01807_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_94_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07345__A3 _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08630_ as2650.stack\[12\]\[3\] _03305_ _03306_ as2650.stack\[13\]\[3\] _03332_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06886__I _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05842_ _00850_ net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05790__I as2650.debug_psl\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_169_Left_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ as2650.stack\[15\]\[1\] _03264_ _03254_ as2650.stack\[14\]\[1\] _03256_ _03265_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_89_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05773_ _00770_ _00783_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07512_ _02320_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08492_ _01274_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_112_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_146_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07443_ _02237_ _02269_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08058__A1 net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07374_ _02191_ _02209_ _02210_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_169_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09113_ _03752_ _03802_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06325_ _01244_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07805__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11032__I _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09044_ _01748_ _03735_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06256_ _01129_ _01224_ _01228_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_130_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06187_ _01159_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10168__A2 _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05965__I _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08230__A1 _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_165_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08781__A2 _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ _01519_ _01465_ _04579_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_141_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09877_ _04525_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08828_ as2650.stack\[11\]\[10\] _03461_ _03514_ as2650.stack\[10\]\[10\] _03523_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06796__I _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_120_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _00641_ _03226_ _01878_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output216_I net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11770_ _00549_ clknet_leaf_3_wb_clk_i as2650.stack\[14\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08717__S _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10721_ as2650.stack\[8\]\[5\] _05197_ _05199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06847__A2 _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08049__A1 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10652_ _04904_ _05146_ _05149_ _04908_ _05151_ _05155_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_TAPCELL_ROW_118_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10583_ as2650.stack\[15\]\[13\] _05106_ _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_114_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06036__I _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07272__A2 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11204_ _05459_ _05562_ _05564_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11135_ _01685_ _05186_ _04522_ _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11108__A1 _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06783__A1 _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11066_ _01958_ _05477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10017_ as2650.stack\[10\]\[0\] _04627_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10919_ _04910_ _05276_ _05356_ _05357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10398__A2 _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06110_ _01082_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_54_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07090_ _01974_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08460__A1 as2650.ivectors_base\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06041_ _01026_ net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_140_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09800_ _04480_ _02620_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_61_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07992_ _02725_ _01791_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_158_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_163_Right_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06943_ _01856_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09731_ _03728_ _04415_ _04281_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08515__A2 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _04339_ _04347_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06874_ _01791_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06526__A1 _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08613_ _02704_ _03108_ _03240_ _03281_ _03315_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05825_ _00830_ _00831_ _00832_ _00833_ _00734_ _00704_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_09593_ _01779_ _01599_ _03633_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_94_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11027__I _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08544_ _02489_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05756_ _00766_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08475_ as2650.ivectors_base\[9\] _03180_ _03182_ _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05687_ _00687_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_110_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07426_ _02078_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_154_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07357_ _02181_ wb_counter\[12\] _02195_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ _01096_ _01159_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07288_ _02114_ _02131_ _02134_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_80_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_80_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_167_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ _03716_ _03718_ _03703_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06239_ _01211_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05695__I _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10561__A2 _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09929_ net140 _01466_ _04572_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08506__A2 _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11753_ _00532_ clknet_leaf_94_wb_clk_i as2650.regs\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10704_ _01694_ _05186_ _01962_ _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_83_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07493__A2 _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11684_ _00468_ clknet_leaf_20_wb_clk_i as2650.stack\[8\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10635_ _02590_ _05141_ _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_36_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10566_ as2650.stack\[15\]\[8\] _05096_ _05097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10497_ _04629_ _05046_ _05050_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08745__A2 _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10016__I _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10552__A2 _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11118_ _05459_ _05508_ _05510_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_53_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__C _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11049_ _01912_ _05465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput7 bus_in_gpios[6] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05610_ as2650.indirect_target\[9\] _00621_ _00623_ as2650.PC\[9\] _00624_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06590_ _01086_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_52_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08260_ _01138_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_47_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08681__B2 as2650.stack\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07211_ net70 _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_rebuffer2_I net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08191_ _01001_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07142_ _02023_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08433__A1 _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07073_ as2650.stack\[11\]\[1\] _01975_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07787__A3 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06995__A1 as2650.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06024_ _00889_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06404__I net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_147_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07975_ _02731_ _02702_ _02732_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_96_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09714_ _04352_ _04398_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06926_ _01838_ _01805_ _01839_ _01840_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_143_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07235__I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06857_ _01718_ _01767_ _01775_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09645_ _04329_ _04330_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ as2650.regs\[2\]\[3\] _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09576_ _04255_ _04261_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06788_ _01262_ _01238_ _01323_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08527_ _03222_ _03225_ _03231_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05739_ _00709_ _00750_ _00751_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_93_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ _03163_ _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07409_ _02081_ wb_counter\[19\] _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ as2650.stack\[0\]\[14\] _02493_ _02500_ as2650.stack\[1\]\[14\] _02506_ _03110_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_163_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_169_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10420_ _04798_ _04799_ _01382_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08424__A1 as2650.stack\[15\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output283_I net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10231__A1 _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10351_ _02626_ _04728_ _04764_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10282_ _04360_ _04806_ _04858_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08727__A2 _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07145__I _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10298__A1 _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11805_ _00584_ clknet_leaf_110_wb_clk_i as2650.stack\[9\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11736_ _00520_ clknet_leaf_23_wb_clk_i as2650.stack\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_139_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11667_ _00451_ clknet_leaf_80_wb_clk_i as2650.regs\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10618_ as2650.stack\[7\]\[9\] _05130_ _05132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08704__I _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11598_ _00382_ clknet_leaf_123_wb_clk_i as2650.stack\[2\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10549_ _01819_ _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_122_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06977__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06729__A1 net250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_119_wb_clk_i_I clknet_4_10__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10525__A2 _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07760_ _02528_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_155_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06711_ _01390_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__10289__A1 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10289__B2 _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07691_ net234 _01628_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09430_ _04100_ _04109_ _04113_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_71_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06642_ _01576_ _01578_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_49_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09361_ _03993_ _03996_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06573_ _01517_ _01522_ _01521_ net156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_47_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08312_ _03021_ _02577_ _03022_ net209 _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_19_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_19_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ _03904_ _03905_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_151_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11581__CLK clknet_leaf_92_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08243_ _02969_ _02628_ _02976_ net200 _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08406__A1 _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08174_ _01167_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11005__A3 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07125_ _02008_ _02012_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07056_ _01712_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_1474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput130 net130 RAM_start_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput141 net141 bus_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput152 net152 bus_data_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06007_ _01007_ net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05640__A1 _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput163 net163 io_oeb[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput174 net174 io_out[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_145_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input42_I io_in[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05973__I _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput185 net300 io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput196 net196 la_data_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07393__A1 net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07958_ _02716_ _02678_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__05943__A2 _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06909_ _01823_ _01805_ _01824_ _01783_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07889_ _02637_ _01708_ _02650_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output129_I net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09628_ _01682_ _03720_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09559_ _03667_ _03773_ _03775_ _03637_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_93_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11521_ _00305_ clknet_leaf_68_wb_clk_i as2650.io_bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_110_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06120__A2 _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05849__I3 _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11452_ _00236_ clknet_leaf_35_wb_clk_i as2650.PC\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__I _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10403_ _01657_ _04858_ _04974_ _04975_ _04746_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_34_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08948__A2 _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11383_ _00009_ clknet_leaf_65_wb_clk_i as2650.cycle\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09070__A1 _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10334_ as2650.regs\[5\]\[4\] _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_91_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10265_ _04231_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10196_ _04773_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11454__CLK clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_89_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07687__A2 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05698__A1 _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11125__I _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07439__A2 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11719_ _00503_ clknet_leaf_82_wb_clk_i as2650.regs\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput10 bus_in_serial_ports[1] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08434__I _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput21 bus_in_sid[4] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07478__C _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput32 bus_in_timers[7] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput43 irqs[0] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput54 ram_bus_in[4] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05870__A1 net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput65 rom_bus_in[7] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput76 net395 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput87 net423 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10746__A2 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_137_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_137_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput98 net357 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08930_ _03619_ _03621_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_110_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ _03372_ _03554_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07812_ _01277_ _01364_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_140_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08792_ as2650.stack\[0\]\[9\] _02492_ _02499_ as2650.stack\[1\]\[9\] _02505_ _03488_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_139_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07743_ _02511_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07674_ _02449_ _02450_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07678__A2 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09413_ _00775_ _00793_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10682__A1 _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06625_ as2650.debug_psl\[5\] _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11035__I _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06556_ _01206_ _01207_ _01510_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09344_ _04026_ _04028_ _04029_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10434__A1 _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09275_ _03950_ _03951_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06487_ _01002_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_35_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07150__I1 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ as2650.instruction_args_latch\[1\] _02950_ _02962_ _02958_ _02963_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05861__A1 _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08157_ _02572_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_133_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07108_ _01959_ _01992_ _01997_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _02839_ _02829_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05613__B2 as2650.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ _01946_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10050_ _01912_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_140_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output246_I net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_127_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07118__A1 wb_feedback_delay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10952_ _01729_ _05386_ _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10883_ net189 _04933_ _05323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06341__A2 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08963__B _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06039__I _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08682__C _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10784__I _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07141__I1 net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11504_ _00288_ clknet_leaf_67_wb_clk_i net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_129_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11435_ _00219_ clknet_4_7__leaf_wb_clk_i as2650.page_reg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09043__A1 _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold50_I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11366_ _00162_ clknet_leaf_69_wb_clk_i net228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05604__A1 as2650.indirect_target\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05604__B2 as2650.PC\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10317_ _04224_ _04861_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11297_ _00093_ clknet_leaf_144_wb_clk_i net294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09085__I _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10248_ _04825_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10179_ _04757_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05758__I2 net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08857__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07333__I _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06332__A2 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06410_ _01372_ _01373_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07390_ _02136_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08592__C _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05930__I2 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06341_ _01293_ _01295_ _01289_ _01309_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_44_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09282__A1 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07132__I1 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06096__A1 net234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10967__A2 _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09060_ _03698_ _03700_ _03713_ _03751_ _01538_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_128_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06272_ _01243_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_60_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06635__A3 _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08011_ as2650.indirect_target\[4\] _02761_ _02762_ _02767_ _02630_ _02768_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_71_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__A1 _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09585__A2 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08793__B1 _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _01488_ _01658_ _04591_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08913_ _01389_ _01211_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09893_ as2650.stack\[5\]\[14\] _04546_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08844_ as2650.stack\[3\]\[11\] _03141_ _03143_ as2650.stack\[2\]\[11\] _03538_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05987_ _00973_ _00939_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08775_ as2650.stack\[12\]\[8\] _02526_ _02529_ as2650.stack\[13\]\[8\] _03472_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07726_ _02494_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08848__B2 _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ net92 _02426_ _02434_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06608_ web_behavior\[0\] _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_94_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07588_ wb_counter\[14\] _02379_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__A1 _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09327_ _00817_ _01494_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06539_ _01497_ net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08074__I _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _03939_ _03942_ _03943_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_output196_I net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07823__A2 _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08209_ as2650.warmup\[0\] as2650.warmup\[1\] _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09189_ _00790_ _00896_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09025__A1 _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11220_ _05477_ _05568_ _05573_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_112_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11151_ _05449_ _05529_ _05531_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_129_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10102_ as2650.stack\[3\]\[11\] _04682_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_129_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11082_ _05479_ _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10033_ _01834_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_125_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08677__C _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06478__B _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10646__A1 _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10646__B2 _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10935_ _05290_ _00801_ _01087_ _05372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_98_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold98_I wbs_adr_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10866_ as2650.chirpchar\[1\] _05267_ _04781_ _05307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08067__A2 _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10797_ as2650.stack\[6\]\[9\] _05244_ _05246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10949__A2 _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10019__I _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_124_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08712__I _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ _00202_ clknet_leaf_86_wb_clk_i as2650.warmup\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09567__A2 _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08775__B1 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11349_ _00145_ clknet_leaf_138_wb_clk_i wb_counter\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06250__A1 _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05910_ as2650.regs\[2\]\[4\] _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06890_ _01806_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06002__A1 _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05841_ _00847_ _00848_ _00849_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06553__A2 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05772_ _00661_ _00778_ _00781_ _00748_ _00782_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08560_ _01690_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07063__I _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07511_ _02319_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10637__A1 _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08491_ _01721_ _03195_ _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07502__A1 net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07442_ net282 _02238_ _02268_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07373_ net271 _02197_ _02188_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11460__D _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06069__A1 net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06324_ _01292_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_21_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _01772_ _03049_ _03765_ _03798_ _03800_ _03801_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
Xclkbuf_leaf_152_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_152_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_169_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07805__A2 net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09043_ _01575_ _02475_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_143_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06255_ _01186_ _01227_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06186_ net63 _01153_ _01158_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__10373__B _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08766__B1 _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_165_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09945_ _02791_ _04578_ _04582_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_121_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09876_ _01869_ _04533_ _04538_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08827_ _03515_ _03518_ _03519_ _03521_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_77_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _02702_ _02830_ _03399_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_1623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output111_I net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07709_ _02477_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_output209_I net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09494__A1 _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08689_ _03324_ _03386_ _03388_ _01445_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_138_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10720_ _05084_ _05196_ _05198_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10651_ as2650.regs\[1\]\[3\] _05155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09246__B2 _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10582_ _01946_ _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09797__A2 _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_75_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09549__A2 _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11203_ as2650.stack\[9\]\[8\] _05563_ _05564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11134_ _05477_ _05514_ _05519_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07980__A1 _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06783__A2 _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11065_ _05475_ _05470_ _05476_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06987__I _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10016_ _04626_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_137_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_4_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__A2 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06299__A1 _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10918_ _05272_ _05354_ _05355_ _05341_ _05356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_54_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07611__I _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10849_ _05284_ _05291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06040_ _01025_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_125_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_100_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07991_ _01453_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_157_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09730_ _04409_ _04414_ _04277_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06942_ _01855_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_78_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09173__B1 _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09661_ _04342_ _04346_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06873_ _01788_ _01790_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__06526__A2 as2650.cycle\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10212__I _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08612_ _01789_ _03283_ _03225_ _03314_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_05824_ _00823_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05734__B1 _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09592_ _04270_ _04276_ _04277_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_19_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08543_ as2650.stack\[3\]\[1\] _03244_ _03246_ as2650.stack\[2\]\[1\] _03247_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05755_ _00765_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05686_ _00699_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08474_ _03174_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_159_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10368__B _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_4_12__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07425_ _02244_ wb_counter\[21\] _02254_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__A1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11043__I _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09779__A2 _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07356_ _02192_ _01780_ _02194_ _02170_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_73_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06307_ _01277_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07287_ _02116_ _02132_ _02133_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_143_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_167_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06238_ _01210_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09026_ _03717_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_167_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08739__B1 _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06169_ _01141_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_125_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output159_I net159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09928_ _04571_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09859_ as2650.stack\[5\]\[0\] _04528_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_1707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_68_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07478__B1 _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11752_ _00531_ clknet_leaf_88_wb_clk_i as2650.chirpchar\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10703_ _01712_ _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10872__I1 _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11683_ _00467_ clknet_leaf_20_wb_clk_i as2650.stack\[8\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10634_ _04698_ _05141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06047__I _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__C _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10565_ _05075_ _05096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_84_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06453__A1 _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10496_ as2650.stack\[1\]\[1\] _05048_ _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06205__A1 net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_109_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06756__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11117_ as2650.stack\[14\]\[8\] _05509_ _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_53_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09093__I _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11048_ _05463_ _05460_ _05464_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput8 bus_in_gpios[7] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10068__A2 _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07469__B1 _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09042__B _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07341__I _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_47_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08681__A2 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07210_ net105 _02006_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08190_ _02866_ _02932_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06692__A1 _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07141_ net100 net134 _02020_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_148_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08433__A2 _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09630__A1 _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06444__A1 _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold102_I wbs_dat_i[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07072_ _01737_ _01973_ _01976_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06023_ _01014_ net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_168_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08197__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06747__A2 _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07944__A1 _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07974_ _02643_ _02730_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09713_ _04338_ _04343_ _04397_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_103_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06925_ _01782_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_143_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_143_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11038__I _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09161__A3 _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09644_ _01560_ _02790_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06856_ _01769_ _01770_ _01774_ _01717_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_155_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05807_ _00816_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ _04256_ _04260_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_102_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06787_ _01253_ _01455_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_17_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_156_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_156_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08526_ _02649_ _03064_ _03228_ _01045_ _03230_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__10059__A2 _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05738_ _00693_ as2650.regs\[7\]\[6\] _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08457_ _01857_ _03164_ _03170_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05669_ _00669_ _00671_ _00673_ _00682_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_149_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07408_ _02084_ net115 _02087_ _01902_ _02146_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_4_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08388_ as2650.stack\[3\]\[14\] _01693_ _01969_ as2650.stack\[2\]\[14\] _03109_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_162_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ net267 _02166_ _02160_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08424__A2 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05869__S0 net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ _01397_ _04791_ _04826_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_143_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output276_I net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06986__A2 _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09009_ _01263_ _02561_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10281_ _04847_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_143_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08188__A1 _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09924__A2 net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07426__I _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09688__A1 _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11804_ _00583_ clknet_leaf_150_wb_clk_i as2650.stack\[9\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11735_ _00519_ clknet_leaf_24_wb_clk_i as2650.stack\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09860__A1 _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06674__A1 net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_148_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11666_ _00450_ clknet_leaf_94_wb_clk_i as2650.regs\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10617_ _05094_ _05129_ _05131_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11597_ _00381_ clknet_leaf_129_wb_clk_i as2650.stack\[2\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10548_ _05082_ _05074_ _05083_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10479_ _05018_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08179__A1 _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_1640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07926__A1 _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06710_ _01626_ _01627_ _01635_ _01636_ net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_07690_ _02459_ _02460_ _02004_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_95_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08351__A1 _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10697__I _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06641_ _01129_ _01276_ _01577_ _01214_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_17_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09360_ _04010_ _04011_ _04045_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06572_ _01523_ net158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_1368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08103__A1 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08311_ _02913_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09291_ _03974_ _03975_ _03976_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_151_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08242_ _02951_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_1655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_59_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_59_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08173_ _01748_ _02914_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09603__A1 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06417__A1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ net66 net67 _02011_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_82_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06968__A2 _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07055_ _01930_ _01959_ _01960_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_149_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput120 net120 RAM_end_addr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_149_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput131 net131 RAM_start_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput142 net142 bus_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06006_ _01006_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07217__I0 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput153 net153 bus_data_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09906__A2 _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput164 net303 io_oeb[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_145_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput175 net175 io_out[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput186 net298 io_out[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput197 net197 la_data_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input35_I io_in[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07957_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_138_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07690__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05794__I3 _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06908_ _01569_ _01809_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07888_ _02638_ _02641_ _02649_ _01320_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09627_ _04295_ _04299_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_168_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06839_ _01718_ _01746_ _01758_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XPHY_EDGE_ROW_90_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09558_ _03637_ _03666_ _04243_ _01231_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_78_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08509_ _02554_ _02555_ _03213_ _01219_ _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_136_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08645__A2 _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09489_ _04035_ _04038_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11520_ _00304_ clknet_leaf_75_wb_clk_i as2650.ext_io_addr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11451_ _00235_ clknet_leaf_32_wb_clk_i as2650.ivectors_base\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10402_ _03745_ _04731_ _04847_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11382_ _00008_ clknet_leaf_66_wb_clk_i as2650.cycle\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09070__A2 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10333_ _04880_ _04789_ _04904_ _04835_ _04908_ _04840_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_TAPCELL_ROW_91_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08540__I _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ as2650.regs\[5\]\[2\] _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_63_1694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08176__A4 _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10195_ _04773_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08333__A1 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10691__A2 _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_44_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08636__A2 _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09833__A1 _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11718_ _00502_ clknet_leaf_80_wb_clk_i as2650.regs\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput11 bus_in_serial_ports[2] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11649_ _00433_ clknet_4_10__leaf_wb_clk_i as2650.stack\[7\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput22 bus_in_sid[5] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput33 io_in[0] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput44 irqs[1] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput55 ram_bus_in[5] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05870__A2 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput66 wb_rst_i net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput77 net397 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput88 net424 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07072__A1 _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput99 net361 net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_161_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05622__A2 _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08860_ _01916_ _01449_ _03483_ _03551_ _03553_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08021__B1 _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07811_ _02579_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_106_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_106_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08791_ as2650.stack\[3\]\[9\] _01692_ _02512_ as2650.stack\[2\]\[9\] _03487_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_97_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ _01965_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__A1 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07673_ net221 _01638_ _01611_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08875__A2 _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09412_ _04097_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06624_ wb_debug_cc _01565_ _01540_ _01566_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_149_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09343_ _01500_ _01495_ _01018_ _04027_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_75_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06555_ _01203_ _01509_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_158_Right_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10434__A2 _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09274_ _03874_ _03883_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_63_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06486_ _01254_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_118_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08225_ _02904_ _02960_ _02961_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08156_ _02632_ _02902_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07107_ as2650.stack\[11\]\[15\] _01993_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08087_ _02800_ _02825_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07038_ _00958_ _01843_ _01945_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_140_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output239_I net239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ _03607_ _03647_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10370__A1 _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07118__A2 _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_123_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_123_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10951_ _03158_ _04432_ _03440_ _04189_ _05386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_138_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06877__A1 _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10882_ _03311_ _05321_ _05322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_168_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_80_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_136_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06629__A1 _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09140__B _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_2__f_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11503_ _00287_ clknet_leaf_59_wb_clk_i as2650.trap vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_53_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_93_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11434_ _00218_ clknet_leaf_56_wb_clk_i as2650.instruction_args_latch\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09043__A2 _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_78_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11365_ _00161_ clknet_leaf_68_wb_clk_i net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_4_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10316_ _01626_ _04848_ _04890_ _04891_ _04746_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_11296_ _00092_ clknet_leaf_144_wb_clk_i net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10305__I _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10247_ _01083_ _04372_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_33_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10178_ _01165_ _02934_ _01795_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10361__A1 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05758__I3 _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08873__C _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09806__A1 _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06340_ _01298_ _01303_ _01306_ _01308_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_57_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05930__I3 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09282__A2 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06271_ _01242_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_72_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08010_ _02766_ _02678_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_147_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09034__A2 _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07045__A1 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09961_ net225 _01545_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _03603_ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_141_1478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10215__I _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09892_ _01947_ _04545_ _04548_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08843_ _03284_ _03535_ _03536_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08774_ as2650.stack\[8\]\[8\] _03249_ _03251_ as2650.stack\[9\]\[8\] _03252_ _03471_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05986_ _00987_ net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07725_ _01873_ as2650.debug_psu\[1\] _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_139_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11046__I _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07656_ wb_counter\[28\] _02436_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_0_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06607_ _01552_ clknet_1_1__leaf__01549_ net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_165_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07587_ _02373_ _02380_ _02381_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06584__B _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05979__I _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09326_ _04009_ _04010_ _04011_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06538_ _01496_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10958__A3 _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ _00792_ _00875_ _03938_ _03892_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06469_ _01427_ _01431_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08208_ as2650.warmup\[0\] _02947_ _01034_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09188_ _03869_ _03873_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA_output189_I net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07036__A1 net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08139_ _02866_ _02887_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_1643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11150_ as2650.stack\[13\]\[4\] _05530_ _05531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05598__A1 _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10101_ _04651_ _04681_ _04685_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_73_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11081_ _05173_ _05480_ _05482_ _05486_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_41_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10032_ _04635_ _04636_ _04638_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_125_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10343__A1 _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09850__S _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06478__C _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10934_ _04959_ _04960_ _05291_ _05371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_131_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10865_ _03268_ _05266_ _05304_ _05305_ _05306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09264__A2 _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10796_ _05094_ _05243_ _05245_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07275__A1 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_10_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07027__A1 _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11417_ _00201_ clknet_leaf_86_wb_clk_i as2650.warmup\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06513__I _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11348_ _00144_ clknet_leaf_138_wb_clk_i wb_counter\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05589__A1 as2650.relative_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11279_ _00075_ clknet_leaf_103_wb_clk_i net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_103_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06002__A2 _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05840_ _00724_ as2650.regs\[6\]\[0\] _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05771_ _00748_ as2650.instruction_args_latch\[6\] _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07510_ net70 _02065_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08490_ _03192_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10637__A2 _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07502__A2 _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07441_ _02239_ _02266_ _02267_ _02094_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_58_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07372_ _02181_ wb_counter\[14\] _02208_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ _03785_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06069__A2 _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06323_ _01041_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_21_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11062__A2 _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _03728_ _03731_ _03733_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06254_ _01226_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_115_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08215__B1 net195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06185_ _01111_ _01157_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_169_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_121_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_121_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09944_ _01520_ _04576_ _04579_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_165_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08518__A1 _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09875_ as2650.stack\[5\]\[7\] _04534_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10325__A1 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08826_ as2650.stack\[4\]\[10\] _03516_ _03517_ as2650.stack\[5\]\[10\] _03520_ _03521_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA_clkbuf_leaf_93_wb_clk_i_I clknet_4_10__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_120_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08757_ _02999_ _03453_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05969_ net226 net245 _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_119_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07708_ _02474_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10628__A2 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08688_ _01831_ _03387_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_68_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09494__A2 _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05703__S _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07639_ _02320_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_1344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08085__I _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10650_ _04874_ _05146_ _05149_ _04879_ _05151_ _05154_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_113_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07257__A1 _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09309_ _03985_ _03893_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10581_ _05104_ _05105_ _05107_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11202_ _05550_ _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11133_ as2650.stack\[14\]\[15\] _05515_ _05519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08509__A1 _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11064_ as2650.stack\[0\]\[14\] _05471_ _05476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10316__A1 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10015_ _04623_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07164__I _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__A3 _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10917_ _04173_ _04963_ _05355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06508__I _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10848_ _03812_ _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07248__A1 _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_138_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10779_ as2650.stack\[6\]\[2\] _05232_ _05235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08748__A1 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07990_ _02718_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06941_ _00727_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__A1 _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09660_ _04343_ _04344_ _04345_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09173__B2 _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06872_ _01719_ _01762_ _01789_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_2_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08920__A1 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ _01275_ _03287_ _03313_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_2_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05823_ net198 _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05734__A1 _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09591_ _03160_ _03768_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05734__B2 _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08542_ _03245_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_49_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05754_ _00764_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_132_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08473_ _00915_ _03179_ _03181_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_158_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05685_ as2650.cycle\[0\] _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_65_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07424_ _02212_ _02252_ _02253_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09228__A2 _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07355_ net125 _02168_ _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06306_ _01205_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07286_ wb_reset_override_en _02124_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09025_ _02579_ _02566_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_167_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06237_ _01115_ _01209_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_167_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input65_I rom_bus_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08739__B2 as2650.stack\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06168_ _01139_ _01140_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07411__A1 net276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06099_ _00999_ _01000_ _01003_ _01075_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_102_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09927_ _01546_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_121_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__A1 _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09858_ _04527_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_107_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output221_I net221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08809_ _01895_ _02723_ _03277_ _03504_ _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_68_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_68_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _01902_ _02617_ _03794_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07478__A1 as2650.wb_hidden_rom_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11751_ _00004_ clknet_leaf_88_wb_clk_i as2650.chirpchar\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07478__B2 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10702_ _05179_ _05184_ _05185_ _00695_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_95_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06150__A1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11682_ _00466_ clknet_leaf_131_wb_clk_i as2650.stack\[8\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11026__A2 _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ _05112_ _05135_ _05140_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10564_ _05073_ _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_134_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06453__A2 _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ _04621_ _05046_ _05049_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11116_ _05496_ _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_21_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05964__A1 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09155__A1 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11047_ as2650.stack\[0\]\[9\] _05461_ _05464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08902__A1 _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput9 bus_in_serial_ports[0] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_95_1365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07622__I _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09702__I0 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06238__I _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06692__A2 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11017__A2 _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07140_ _02022_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10776__A1 _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07071_ as2650.stack\[11\]\[0\] _01975_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06022_ _01013_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_51_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_147_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07973_ _02726_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09712_ _04339_ _04342_ _04345_ _04396_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_06924_ _01560_ _01809_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_143_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09643_ _03159_ _02802_ _03707_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_39_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06855_ _01772_ _01773_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06857__B _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05806_ _00815_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_74_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _04257_ _04258_ _04259_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06786_ _01706_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_102_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08525_ _03229_ _02711_ _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_156_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05737_ as2650.regs\[3\]\[6\] _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_72_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08456_ as2650.ivectors_base\[3\] _03165_ _03167_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05668_ net38 _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08564__S _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07180__I0 net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07407_ _02066_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11008__A2 _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08387_ _03063_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05599_ _00605_ _00608_ _00609_ _00612_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_45_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07338_ _02155_ wb_counter\[10\] _02178_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ _02010_ _02086_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__S1 _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09008_ _03699_ _02924_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_63_1832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10280_ _04849_ _04852_ _04856_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output171_I net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08188__A2 _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05936__B _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09688__A2 _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _00582_ clknet_leaf_150_wb_clk_i as2650.stack\[9\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08112__A2 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11734_ _00518_ clknet_leaf_7_wb_clk_i as2650.stack\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07171__I0 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11665_ _00449_ clknet_leaf_99_wb_clk_i as2650.regs\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10616_ as2650.stack\[7\]\[8\] _05130_ _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11596_ _00380_ clknet_leaf_128_wb_clk_i as2650.stack\[2\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07623__A1 net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10547_ as2650.stack\[15\]\[3\] _05076_ _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08820__B1 _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10478_ _04653_ _05032_ _05037_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_55_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08179__A2 _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05937__A1 _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10930__A1 _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11139__I _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10043__I _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08876__C _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06640_ _01224_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_2_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07352__I _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06571_ as2650.io_bus_we _01522_ _01521_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_08310_ _03033_ _03035_ _03028_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09290_ _03959_ _03960_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_118_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_151_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _01485_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08183__I as2650.instruction_args_latch\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08172_ _01249_ _01242_ _02914_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07123_ _02009_ _02010_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05625__B1 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07054_ as2650.stack\[12\]\[15\] _01941_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_99_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_149_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput110 net110 RAM_end_addr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_105_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_149_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput121 net121 RAM_end_addr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_3_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06005_ _01005_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput132 net132 RAM_start_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput143 net143 bus_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_144_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07217__I1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_28_wb_clk_i clknet_4_6__leaf_wb_clk_i clknet_leaf_28_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput154 net154 bus_data_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput165 net165 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput176 net176 io_out[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput187 net187 io_out[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput198 net198 la_data_out[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__11049__I _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A1 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07956_ _02714_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input28_I bus_in_timers[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06907_ _00803_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07887_ _02644_ _02646_ _02648_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08878__B1 _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06838_ _01747_ _01753_ _01757_ _01734_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_09626_ _04309_ _04311_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ _01282_ _03638_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06769_ _01689_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08508_ _03206_ _03212_ _02549_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09488_ _04039_ _04040_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_52_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08439_ as2650.insin\[7\] _02612_ _02463_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07853__A1 _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11450_ _00234_ clknet_leaf_31_wb_clk_i as2650.ivectors_base\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_134_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10401_ _04849_ _04970_ _04973_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11381_ _00005_ clknet_leaf_65_wb_clk_i as2650.cycle\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10332_ _04906_ _04907_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07865__C _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10263_ _00863_ _04789_ _04834_ _04835_ _04839_ _04840_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_79_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10194_ _04772_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09530__A1 _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08268__I _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09601__B _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11717_ _00501_ clknet_leaf_78_wb_clk_i as2650.regs\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06516__I as2650.cycle\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11648_ _00432_ clknet_leaf_89_wb_clk_i as2650.stack\[7\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput12 bus_in_serial_ports[3] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput23 bus_in_sid[6] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput34 io_in[10] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09597__A1 _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput45 irqs[2] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11579_ _00363_ clknet_leaf_80_wb_clk_i as2650.regs\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput56 ram_bus_in[6] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput67 net408 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_64_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput78 net401 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput89 net421 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08731__I _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09048__B _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__A1 as2650.stack\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07347__I _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06251__I _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09364__A4 _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10364__C1 _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07810_ _02578_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08572__A2 _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08790_ _01895_ _03485_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_140_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07741_ _02509_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07672_ _01538_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09521__B2 _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_146_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_146_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10131__A2 _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09411_ _03922_ _04095_ _04096_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06623_ as2650.insin\[6\] wb_debug_cc _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _01496_ _01018_ _04027_ _01500_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06554_ _00688_ _01228_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_158_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09824__A2 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06638__A2 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09273_ _03952_ _03957_ _03958_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06485_ _01335_ _01447_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ as2650.instruction_args_latch\[1\] _02955_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09588__A1 _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08155_ _02900_ _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07106_ _01954_ _01992_ _01996_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08086_ _02827_ _01892_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_67_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07037_ _01943_ _01770_ _01944_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_100_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08012__A1 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06574__A1 as2650.io_bus_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _03677_ _03678_ _03679_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10370__A2 _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output134_I net134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_127_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07939_ _01334_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08315__A2 _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ _05295_ _05376_ _05385_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_123_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09609_ as2650.debug_psu\[7\] _02465_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06877__A2 _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10881_ _05265_ _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08079__A1 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08079__B2 as2650.indirect_target\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_136_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09815__A2 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07826__A1 _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11502_ _00286_ clknet_leaf_117_wb_clk_i as2650.stack\[5\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09848__S _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__A1 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11433_ _00217_ clknet_leaf_56_wb_clk_i as2650.instruction_args_latch\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11364_ _00160_ clknet_leaf_141_wb_clk_i wb_counter\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10315_ _03858_ _04806_ _04858_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11295_ _00091_ clknet_leaf_144_wb_clk_i net292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10246_ _04791_ _04823_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10177_ _04719_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_33_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07116__B _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06317__A1 _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10113__A2 _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06270_ _00969_ _00998_ _01075_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_127_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08793__A2 _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09960_ _01649_ _04590_ _01088_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_1570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08911_ _03600_ _03602_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_0_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09891_ as2650.stack\[5\]\[13\] _04546_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09742__A1 _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08842_ _01917_ _03512_ _01916_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_83_wb_clk_i_I clknet_4_15__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08773_ as2650.stack\[11\]\[8\] _03466_ _03462_ as2650.stack\[10\]\[8\] _03470_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05985_ _00981_ _00985_ _00986_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07724_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07655_ wb_counter\[26\] wb_counter\[27\] _02429_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06606_ _01551_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07586_ net398 _02376_ _02368_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07540__I _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09325_ _01014_ _01015_ _01494_ _01489_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_36_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06537_ _01495_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06156__I _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09256_ _03930_ _03940_ _03941_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08481__A1 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06468_ _01428_ _01430_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08207_ as2650.warmup\[1\] _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_43_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09187_ _03872_ _03870_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08608__I0 _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06399_ _01141_ _01150_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_116_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08138_ as2650.ivectors_base\[8\] _02852_ _02886_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_47_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10040__A1 as2650.stack\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08069_ as2650.indirect_target\[7\] _02654_ _02657_ _02815_ _02822_ _02823_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_31_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10100_ as2650.stack\[3\]\[10\] _04682_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_73_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_73_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output251_I net251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11080_ as2650.regs\[7\]\[3\] _05486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_129_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10031_ as2650.stack\[10\]\[4\] _04637_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09733__A1 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05770__A2 _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10933_ as2650.regs\[4\]\[5\] _05288_ _05370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08546__I _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10864_ _01351_ _05265_ _05305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_wire300_I net185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10795_ as2650.stack\[6\]\[8\] _05244_ _05245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_26_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_128_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07275__A2 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08472__A1 as2650.ivectors_base\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08281__I _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11416_ _00200_ clknet_leaf_87_wb_clk_i net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_39_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10031__A1 as2650.stack\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11347_ _00143_ clknet_leaf_107_wb_clk_i wb_counter\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08775__A2 _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11278_ _00074_ clknet_leaf_103_wb_clk_i net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10229_ _04794_ _04802_ _04805_ _04806_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_20_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05770_ _00780_ _00618_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05761__A2 net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07440_ _02081_ wb_counter\[24\] _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06710__A1 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_138_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ _02174_ _02206_ _02207_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_73_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09110_ _03769_ _03799_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06322_ _01291_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ _03732_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10270__A1 _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06253_ _01225_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08405__B _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08191__I _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08215__A1 _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06184_ net34 _01154_ _01156_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_130_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09963__A1 net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08766__A2 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_147_Left_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09943_ _02781_ _04578_ _04581_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08518__A2 _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09874_ _01853_ _04533_ _04537_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08825_ _02518_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__11057__I _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05968_ _00971_ net245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08756_ _03068_ _03095_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input10_I bus_in_serial_ports[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08794__C _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07707_ _01576_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05899_ _00904_ _00900_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_55_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08687_ _01813_ _03363_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_156_Left_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09494__A3 _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07638_ _02407_ _02421_ _02422_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07569_ wb_counter\[11\] _02364_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_118_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09308_ _03931_ _00897_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_118_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07257__A2 net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10580_ as2650.stack\[15\]\[12\] _05106_ _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _03916_ _03924_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_88_1598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08206__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06614__I _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11201_ _05548_ _05562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_165_Left_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11132_ _05475_ _05514_ _05518_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08509__A2 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05674__B _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11063_ _01953_ _05475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08050__B _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__B1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10014_ _04624_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08276__I _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10916_ _05351_ _05352_ _05353_ _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08693__A1 _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10847_ as2650.regs\[4\]\[0\] _05288_ _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_1478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07248__A2 net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08445__A1 _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10778_ _05078_ _05230_ _05234_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__A2 _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09945__A1 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08748__A2 _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06759__A1 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10555__A2 _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06940_ _01803_ _01853_ _01854_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09056__B _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I bus_in_gpios[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06871_ as2650.PC\[2\] _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_2_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05822_ _00817_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_08610_ _01765_ _03288_ _03311_ _03312_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09590_ _04272_ _04275_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05734__A2 _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08541_ _01965_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05753_ _00691_ as2650.regs\[4\]\[6\] _00763_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_136_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08472_ as2650.ivectors_base\[8\] _03180_ _03175_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05684_ _00688_ _00697_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07090__I _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_158_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07423_ _02124_ _01931_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07354_ _02120_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_18_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_154_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08436__A1 as2650.insin\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__B _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06305_ _00680_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07285_ net132 _02119_ _02122_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09024_ _03715_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06236_ _01095_ _01122_ _01123_ _01126_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_115_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08739__A2 _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06167_ as2650.insin\[7\] _01096_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input58_I rom_bus_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06098_ _01074_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_22_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09926_ _01465_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_102_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__A2 _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09857_ _04524_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_107_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_4_14__f_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08808_ _03483_ _03501_ _03503_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_107_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__A2 _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09788_ _04463_ _04469_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_68_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output214_I net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08739_ as2650.stack\[12\]\[7\] _02489_ _02496_ as2650.stack\[13\]\[7\] _03437_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_64_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08096__I _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11750_ _00003_ clknet_leaf_88_wb_clk_i as2650.chirpchar\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10701_ _05178_ _05184_ _05185_ _00750_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_90_1499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11681_ _00465_ clknet_leaf_33_wb_clk_i as2650.stack\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10632_ as2650.stack\[7\]\[15\] _05136_ _05140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08427__A1 _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07868__C _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10234__A1 _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08978__A2 _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10563_ _01882_ _05094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_wire298_I net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06453__A3 _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10494_ as2650.stack\[1\]\[0\] _05048_ _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11115_ _05494_ _05508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05964__A2 net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11046_ _01898_ _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08902__A2 _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_1518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09702__I1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06141__A2 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ _01974_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_113_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06021_ _00816_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10528__A2 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_147_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07972_ _02726_ _01791_ _02729_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_09711_ _02658_ _01608_ _01621_ _02676_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06923_ _01837_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_103_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09642_ _03717_ _04327_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06854_ _01751_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05805_ as2650.regs\[1\]\[3\] as2650.regs\[5\]\[3\] _00800_ _00815_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06785_ _01250_ _01702_ _01705_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09573_ net210 _01625_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_102_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05736_ _00659_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08524_ _00641_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_156_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08657__B2 as2650.stack\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05667_ net58 _00666_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_4
X_08455_ _01838_ _03164_ _03169_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07180__I1 net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07406_ _02077_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08386_ _02702_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_110_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05598_ _00610_ _00593_ _00596_ _00603_ _00611_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_110_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10395__B _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07337_ _02174_ _02176_ _02177_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_151_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _02115_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_60_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06219_ _01103_ _01180_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09007_ _02587_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07199_ _02055_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07196__S _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05946__A2 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09909_ _04556_ net149 _04557_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05952__B as2650.instruction_args_latch\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07699__A2 _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08819__I _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i clknet_4_9__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10289__C _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11802_ _00581_ clknet_leaf_150_wb_clk_i as2650.stack\[9\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08648__A1 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09696__I0 net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11733_ _00517_ clknet_leaf_7_wb_clk_i as2650.stack\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07320__A1 net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07171__I1 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11664_ _00448_ clknet_leaf_99_wb_clk_i as2650.regs\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07871__A2 _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10615_ _05117_ _05130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11595_ _00379_ clknet_4_3__leaf_wb_clk_i as2650.stack\[2\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold66_I wbs_adr_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10546_ _01800_ _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10477_ as2650.stack\[2\]\[11\] _05033_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_55_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11183__A2 _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11029_ _05440_ _05451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08887__A1 _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06362__A2 _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06570_ _01519_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_73_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08240_ _02623_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_111_1635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_1657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05873__A1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08171_ _01998_ as2650.indexed_cyc\[0\] _02915_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_12_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07122_ net68 _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__B2 _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _01958_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_1553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput111 net111 RAM_end_addr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06004_ _00999_ _01004_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xoutput122 net122 RAM_start_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07808__I _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput133 net133 RAM_start_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput144 net144 bus_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput155 net155 bus_we_gpios vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07378__A1 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput166 net166 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput177 net177 io_out[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput188 net188 la_data_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_103_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput199 net199 la_data_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06050__A1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A2 _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_68_wb_clk_i clknet_4_13__leaf_wb_clk_i clknet_leaf_68_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07955_ _01110_ _01112_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_157_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06906_ _01803_ _01820_ _01822_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07886_ _02639_ _02647_ _02602_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09625_ _01923_ _02466_ _02619_ _04310_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_116_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06837_ _01755_ _01756_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07550__A1 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09556_ _03822_ _03829_ _04241_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06768_ _01688_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10437__A1 _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08507_ _03207_ _03208_ _03209_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05719_ _00679_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_52_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06699_ _01625_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_17_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09487_ _04043_ _04172_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08438_ _02992_ _01337_ _03152_ _03153_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_138_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08369_ _01147_ _03069_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10400_ _04853_ _04972_ _04742_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11380_ _00176_ clknet_leaf_47_wb_clk_i as2650.indirect_target\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output281_I net281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09850__I0 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10331_ _04160_ _04783_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_91_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10262_ _04770_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06622__I _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07369__A1 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ _01727_ _01750_ _03735_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_44_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08318__B1 _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06592__A2 as2650.cycle\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08869__A1 _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07541__A1 net362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08097__A2 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11716_ _00500_ clknet_leaf_80_wb_clk_i as2650.regs\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11647_ _00431_ clknet_leaf_89_wb_clk_i as2650.stack\[7\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput13 bus_in_serial_ports[4] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_37_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput24 bus_in_sid[7] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09597__A2 _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput35 io_in[11] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput46 irqs[3] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11578_ _00362_ clknet_leaf_92_wb_clk_i as2650.regs\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput57 ram_bus_in[7] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput68 net410 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput79 net385 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10529_ _04661_ _05065_ _05069_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06532__I _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10364__B1 _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10903__A2 _05339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08887__C _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_4_15__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06583__A2 _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07740_ _02508_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08459__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07363__I _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10667__A1 _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ _02332_ _02447_ _02448_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_36_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10131__A3 _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09410_ _00719_ _00757_ _01030_ _00827_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_88_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06622_ _01564_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_59_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10419__A1 _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06553_ _01203_ _01300_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_48_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _01020_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06484_ _01336_ _01337_ _01446_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09272_ _03945_ _03948_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06638__A3 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_115_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_115_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08223_ _01252_ _02608_ net196 _02952_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08154_ _01949_ _02748_ _02001_ _02794_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09588__A2 _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08796__B1 _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07105_ as2650.stack\[11\]\[14\] _01993_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08085_ _02689_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_67_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_1549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07036_ net192 _01773_ _01782_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06442__I _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input40_I io_in[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08797__C _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08987_ _03610_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06574__A2 _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07938_ _02674_ _02691_ _02697_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_127_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_127_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07869_ _02624_ _02631_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_123_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output127_I net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09608_ as2650.debug_psu\[5\] as2650.debug_psu\[4\] net306 _02546_ _04294_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XTAP_TAPCELL_ROW_84_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10880_ _05262_ _05320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09539_ _03672_ _03668_ _03669_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08079__A2 _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09815__A3 _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06617__I wb_debug_cc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_118_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_136_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11501_ _00285_ clknet_leaf_120_wb_clk_i as2650.stack\[5\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_97_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09928__I _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11432_ _00216_ clknet_leaf_55_wb_clk_i as2650.instruction_args_latch\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09579__A2 _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11363_ _00159_ clknet_leaf_106_wb_clk_i wb_counter\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06262__A1 _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10314_ _04849_ _04886_ _04889_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11294_ _00090_ clknet_leaf_144_wb_clk_i net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10245_ _01616_ _04818_ _04822_ _04815_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_37_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09200__A1 _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10346__B1 _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ _03741_ _04754_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_33_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10897__A1 _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08500__C _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_157_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06317__A2 _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06527__I _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05828__A1 net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09019__A1 _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_1382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07358__I _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08910_ _00803_ _03589_ _03601_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_141_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09890_ _01940_ _04545_ _04547_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09742__A2 _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08841_ _01917_ _01916_ _03512_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_100_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10512__I _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07307__B _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08772_ _03463_ _03465_ _03467_ _03468_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05984_ _00982_ _00983_ _00975_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_154_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07723_ _02491_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06308__A2 _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07505__A1 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ _02423_ _02433_ _02435_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_0_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_0_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06605_ _01550_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07585_ wb_counter\[14\] _02379_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_113_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _00826_ _01016_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_36_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06536_ _01494_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09255_ _03871_ _00897_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06467_ as2650.debug_psl\[7\] _01429_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08481__A2 net204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08206_ _02866_ _02946_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06398_ _01343_ _01362_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_09186_ _01027_ _03871_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08137_ _02837_ _02883_ _02884_ _02885_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_116_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07268__I _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_15__leaf_wb_clk_i clknet_leaf_83_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08068_ _01335_ _02821_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__A1 _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07019_ as2650.stack\[12\]\[11\] _01884_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_12_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_12_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_73_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10030_ _04626_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_105_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output244_I net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09733__A2 _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10932_ _05263_ _05367_ _05368_ _05369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_54_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07731__I _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09249__A1 _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10863_ _05270_ _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10794_ _05231_ _05244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_137_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_101_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06791__B _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11415_ _00199_ clknet_leaf_65_wb_clk_i as2650.extend vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06235__A1 _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11346_ _00142_ clknet_leaf_138_wb_clk_i wb_counter\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09972__A2 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11277_ _00073_ clknet_leaf_112_wb_clk_i net119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_123_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06810__I _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ _04730_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10159_ _04736_ _04737_ _01412_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08160__A1 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07370_ _02183_ _01570_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06321_ as2650.cycle\[5\] _01290_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_31_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06252_ _01210_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09040_ _01779_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_154_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold118_I wbs_dat_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06183_ _01155_ _01154_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08215__A2 _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__A1 _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_169_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09942_ net145 _04576_ _04579_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_165_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09873_ as2650.stack\[5\]\[6\] _04534_ _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08824_ as2650.stack\[7\]\[10\] _03461_ _03462_ as2650.stack\[6\]\[10\] _03519_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08755_ _02674_ _03450_ _03452_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05967_ _00656_ _00970_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_120_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07706_ _01429_ _01224_ _01213_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_90_1615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_130_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_130_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08686_ _03380_ _03385_ _02550_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_94_1795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05898_ _00742_ as2650.instruction_args_latch\[2\] _00859_ _00899_ _00903_ _00904_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__08151__A1 _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07637_ net88 _02410_ _02418_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_66_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07568_ _02358_ _02365_ net374 _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _00792_ _00856_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_76_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06519_ _01117_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_119_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_118_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07499_ wb_reset_override _02305_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09238_ _03919_ _03923_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_79_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output194_I net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09169_ _03855_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_75_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11200_ _05457_ _05556_ _05561_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11210__A1 _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09954__A2 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11131_ as2650.stack\[14\]\[14\] _05515_ _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07726__I _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09706__A2 _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08509__A3 _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06630__I _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _05473_ _05470_ _05474_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10013_ _04623_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10152__I _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__A1 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10915_ as2650.chirpchar\[4\] _05256_ _05353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08693__A2 _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold96_I wbs_dat_i[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _05287_ _05288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_15_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10777_ as2650.stack\[6\]\[1\] _05232_ _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08445__A2 _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07410__B _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10252__A2 _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10004__A2 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11329_ net364 clknet_leaf_146_wb_clk_i wb_reset_override vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07708__A1 _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11158__I _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06870_ as2650.PC\[3\] _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_160_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05821_ _00814_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08540_ _03210_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05752_ _00690_ _00762_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08133__A1 _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08471_ _03162_ _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_1622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05683_ _00694_ _00695_ _00696_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_72_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08684__A2 _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07422_ net117 _02149_ _02213_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09228__A4 _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07353_ _02009_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09633__A1 _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06304_ _01274_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10243__A2 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07284_ wb_counter\[4\] _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_85_1739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09023_ _01232_ _01512_ _02582_ _02584_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__10237__I _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06235_ _01204_ _01191_ _01206_ _01207_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_131_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_167_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05670__A2 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06166_ _00664_ _01138_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_1463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06097_ _01039_ _01072_ _01073_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_70_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09925_ _01477_ _04428_ _04569_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_121_1659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09856_ _04525_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08372__A1 _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ _03502_ _01893_ _02842_ _03052_ _03241_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_107_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i clknet_4_8__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09787_ net210 _04449_ _04468_ _02598_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_68_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06999_ _01905_ _01786_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ as2650.stack\[8\]\[7\] _03411_ _03412_ as2650.stack\[9\]\[7\] _02502_ _03436_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_96_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08669_ _03074_ _03085_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output207_I net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10700_ _05177_ _05184_ _05185_ _00785_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_152_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10482__A2 _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11680_ _00464_ clknet_leaf_24_wb_clk_i as2650.stack\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10631_ _05110_ _05135_ _05139_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09624__A1 _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _05092_ _05085_ _05093_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10147__I _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10493_ _05047_ _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06453__A4 _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07938__A1 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_15_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11114_ _05457_ _05502_ _05507_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11045_ _05459_ _05460_ _05462_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07191__I _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08115__A1 _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09702__I2 net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08666__A2 _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06141__A3 _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10829_ _05270_ _05271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09615__A1 _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06429__A1 _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10225__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09091__A2 _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10057__I _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06020_ _01012_ net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09918__A2 net152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07929__A1 _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_162_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07971_ _02727_ _02700_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_147_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09710_ _04395_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06922_ _01667_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08354__A1 _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _04303_ _04312_ _04317_ _04326_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_06853_ _01771_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05804_ _00708_ _00812_ _00813_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09572_ _01497_ _01353_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06784_ _01171_ _01704_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_116_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08523_ _03227_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_102_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05735_ _00743_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_77_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07865__B1 _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08454_ as2650.ivectors_base\[2\] _03165_ _03167_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05666_ _00664_ _00678_ _00679_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_65_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07405_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09606__A1 _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08385_ _01102_ _03059_ _01949_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05597_ as2650.indirect_target\[2\] _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_162_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07336_ _02083_ _01755_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10216__A2 _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09082__A2 _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07093__A1 as2650.stack\[11\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07267_ _02112_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_61_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09756__I _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09006_ _03580_ _02919_ _03656_ _03697_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__09909__A2 net149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06218_ _01190_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_104_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07198_ net96 net112 _02051_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06149_ _01118_ _01121_ _01079_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_93_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09908_ _04555_ _01616_ _04559_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09839_ _04515_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11801_ _00580_ clknet_leaf_150_wb_clk_i as2650.stack\[9\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_139_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08648__A2 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09696__I1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11732_ _00516_ clknet_leaf_4_wb_clk_i as2650.stack\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07856__B1 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07320__A2 _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11663_ _00447_ clknet_leaf_97_wb_clk_i as2650.regs\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_153_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08056__B _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10614_ _05115_ _05129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11594_ _00378_ clknet_leaf_128_wb_clk_i as2650.stack\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _05080_ _05074_ _05081_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08820__A2 _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06831__A1 _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10476_ _04651_ _05032_ _05036_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_55_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10605__I _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07387__A2 _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__A1 _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_4_13__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10391__A1 _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07914__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11028_ _05438_ _05450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10143__A1 _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09300__A3 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05873__A2 _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08170_ _02713_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07121_ net69 _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold100_I wbs_dat_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05625__A2 _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07052_ as2650.page_reg\[2\] _01718_ _01957_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_45_1520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06003_ _01000_ _01003_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput112 net112 RAM_end_addr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_149_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput123 net123 RAM_start_addr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_149_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput134 net134 RAM_start_addr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput145 net145 bus_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput156 net156 bus_we_serial_ports vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_122_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08575__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput167 net167 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_45_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput178 net178 io_out[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput189 net189 la_data_out[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_103_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06050__A2 _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07954_ _02712_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_50_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06905_ as2650.stack\[12\]\[4\] _01821_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07885_ _02643_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10134__A1 _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08878__A2 _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09624_ _03732_ _04307_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_93_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06836_ _01751_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_168_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09555_ _03667_ _03664_ _03665_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_56_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06767_ _01687_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_leaf_37_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_37_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08506_ as2650.stack\[15\]\[0\] _03210_ _02540_ as2650.stack\[14\]\[0\] _03204_ _03211_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05718_ _00705_ _00730_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_108_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09486_ _04032_ _04041_ _04042_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_06698_ _01405_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08437_ _03154_ _03155_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05649_ as2650.cycle\[0\] _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_65_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08368_ _03073_ _03087_ _03089_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_163_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07319_ _02079_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_134_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08299_ _01449_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_95_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05616__A2 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10330_ _04194_ _04774_ _04905_ _04876_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06903__I _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10261_ _04837_ _04838_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_131_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08566__A1 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10192_ _04770_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10373__A1 _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08318__A1 _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_147_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_48_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_48_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09818__A1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11715_ _00499_ clknet_leaf_77_wb_clk_i as2650.regs\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11646_ _00430_ clknet_leaf_124_wb_clk_i as2650.stack\[7\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09046__A2 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 bus_in_serial_ports[5] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_92_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput25 bus_in_timers[0] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput36 io_in[12] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11577_ _00361_ clknet_leaf_89_wb_clk_i as2650.stack\[3\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput47 irqs[4] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__B _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput58 rom_bus_in[0] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07909__I _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput69 net406 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10528_ as2650.stack\[1\]\[14\] _05066_ _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06813__I _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10335__I _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10459_ _05018_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06407__I1 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05873__B _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_140_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07670_ net96 _02340_ _02074_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06621_ as2650.debug_psl\[7\] _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_88_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09340_ _01015_ _01490_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06552_ _01266_ _01506_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06099__A2 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _03945_ _03948_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06483_ _01222_ _01445_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08222_ _02949_ _02959_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_8_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08153_ as2650.indirect_target\[14\] _02757_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_155_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_155_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08796__A1 as2650.stack\[11\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07104_ _01947_ _01992_ _01995_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06723__I _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08084_ _02835_ _02836_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_1528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07035_ _01092_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_12_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10355__A1 _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _03613_ _03642_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input33_I io_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _02692_ _02696_ as2650.irqs_latch\[7\] _01450_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_127_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_127_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07868_ as2650.insin\[5\] _02596_ _02577_ _02600_ _02630_ _02631_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_123_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08720__A1 _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06819_ as2650.stack\[12\]\[0\] _01739_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09607_ _04286_ _04290_ _04291_ _04292_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_84_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07799_ _02567_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_151_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09538_ _01168_ _04218_ _04223_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_66_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09469_ _04153_ _04154_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11500_ _00284_ clknet_leaf_118_wb_clk_i as2650.stack\[5\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11431_ _00215_ clknet_leaf_55_wb_clk_i as2650.instruction_args_latch\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_168_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08787__A1 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11362_ _00158_ clknet_leaf_106_wb_clk_i wb_counter\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06633__I _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10313_ _04853_ _04888_ _04742_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10155__I _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11293_ _00089_ clknet_leaf_155_wb_clk_i net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10244_ _04819_ _04821_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10346__A1 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09200__A2 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10175_ _02922_ _04753_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_98_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08509__B _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06808__I _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05828__A2 _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09019__A2 _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11629_ _00413_ clknet_leaf_21_wb_clk_i as2650.stack\[15\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07639__I _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_1826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07450__A1 net283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10337__A1 _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08840_ _03235_ _03508_ _03533_ _03534_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_110_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06556__A3 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08771_ as2650.stack\[4\]\[8\] _03261_ _03262_ as2650.stack\[5\]\[8\] _03256_ _03468_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05983_ _00982_ _00983_ _00984_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_40_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07722_ _02490_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_75_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09803__B _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07505__A2 _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07653_ net91 _02426_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_1365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06604_ _01076_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07584_ _02378_ _02374_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_152_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09323_ _01029_ _01019_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06535_ _01493_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11065__A2 _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09254_ _00824_ _00815_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10812__A2 _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06466_ _01186_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_145_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08205_ net213 _02945_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09185_ _00912_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_90_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06397_ _01344_ _01361_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08136_ as2650.indirect_target\[12\] _01330_ _02848_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_116_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10576__A1 _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08067_ _02736_ _01456_ _02820_ _02724_ as2650.indirect_target\[7\] _02821_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_77_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07992__A2 _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07018_ _01927_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_73_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_73_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_129_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08601__C _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10703__I _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06547__A3 _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output237_I net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_52_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_52_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08969_ _02601_ _01373_ _01226_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_86_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09497__A2 _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10931_ _04306_ _04308_ _05280_ _05368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_19_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08329__B _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10862_ _05275_ _05303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09249__A2 _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10793_ _05229_ _05243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_149_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09939__I _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06483__A2 _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11414_ _00198_ clknet_leaf_51_wb_clk_i as2650.indirect_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_10_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06235__A2 _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11345_ _00141_ clknet_leaf_141_wb_clk_i wb_counter\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10319__A1 _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11276_ _00072_ clknet_leaf_112_wb_clk_i net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__05994__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10227_ _04803_ _04804_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_105_1590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08932__A1 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10158_ _04703_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10089_ _04639_ _04675_ _04678_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08160__A2 _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06538__I _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06171__A1 _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06320_ _01289_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08999__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06251_ _00688_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07671__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ net55 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_52_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06226__A2 _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A1 _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09941_ _02766_ _04578_ _04580_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_165_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09176__A1 _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10523__I _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _01835_ _04533_ _04536_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08923__A1 _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ as2650.stack\[0\]\[10\] _03516_ _03517_ as2650.stack\[1\]\[10\] _03464_ _03518_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i clknet_4_7__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08754_ _03095_ _03451_ _02667_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_05966_ _00747_ net429 _00955_ _00965_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_120_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07705_ _01130_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_139_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08685_ _03381_ _03382_ _03383_ _03384_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05897_ _00901_ _00902_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07636_ wb_counter\[24\] _02420_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06162__A1 _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07567_ net373 _02361_ _02351_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09306_ _03982_ _03989_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__09100__A1 _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09759__I _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06518_ as2650.cycle\[11\] _01245_ _01478_ _01463_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_118_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07498_ _02310_ net359 _02309_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09237_ _03920_ _03921_ _03922_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_TAPCELL_ROW_79_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06449_ _01411_ _01365_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07662__A1 net392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06465__A2 _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09168_ _01419_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_75_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output187_I net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08119_ _02868_ _02858_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09708__B _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09099_ _01434_ _03786_ _03787_ _03788_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_114_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11130_ _05473_ _05514_ _05517_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09167__A1 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11061_ as2650.stack\[0\]\[13\] _05471_ _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_79_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09706__A3 _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08914__A1 _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A2 _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _01961_ _01962_ _04622_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_4_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07742__I _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08678__B1 _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__A2 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10914_ net191 _04772_ _05270_ _05352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10845_ _03812_ _05285_ _05286_ _05287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_41_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold89_I wbs_dat_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10776_ _05071_ _05230_ _05233_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10788__A1 _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08506__C _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07653__A1 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07410__C _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07917__I _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11328_ net360 clknet_leaf_145_wb_clk_i wb_reset_override_en vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_97_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05967__A1 _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11259_ _00055_ clknet_leaf_150_wb_clk_i net133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_24_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10712__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05820_ _00811_ as2650.instruction_args_latch\[3\] _00749_ _00828_ _00829_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__07652__I _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_167_Right_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05751_ as2650.regs\[0\]\[6\] _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08470_ _03163_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05682_ _00694_ as2650.regs\[7\]\[7\] _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07192__I0 net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07421_ _02190_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_158_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_158_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07352_ _02190_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09633__A2 _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06303_ _01100_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06447__A2 _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07644__A1 _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ _02079_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_155_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07099__I _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09022_ _01221_ _02598_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06234_ _01196_ _01164_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_113_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__A1 _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06165_ _01080_ _01136_ _01137_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__05670__A3 _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07827__I _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06096_ net234 _01038_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__05958__A1 _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09924_ _01313_ net146 as2650.cycle\[7\] _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09855_ _04524_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08806_ _03226_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_107_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06998_ _01908_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_107_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _02521_ _04464_ _04467_ _02484_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05949_ _00745_ as2650.instruction_args_latch\[10\] _00951_ _00953_ _00954_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08737_ as2650.stack\[11\]\[7\] _03428_ _03429_ as2650.stack\[10\]\[7\] _03435_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_154_1458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08124__A2 _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08668_ _01469_ _03350_ _03368_ _03277_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07183__I0 net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07619_ _02357_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_165_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08599_ _02490_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_95_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10630_ as2650.stack\[7\]\[14\] _05136_ _05139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09624__A2 _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10561_ as2650.stack\[15\]\[7\] _05086_ _05093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10492_ _05044_ _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_122_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__I _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05949__A1 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09157__C _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10942__A1 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ as2650.stack\[14\]\[7\] _05503_ _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10163__I _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11044_ as2650.stack\[0\]\[8\] _05461_ _05462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06126__A1 _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07174__I0 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06816__I _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10828_ _04187_ _01729_ _05270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08823__B1 _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10225__A3 _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10759_ _05173_ _05215_ _05217_ _05221_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_82_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_92_wb_clk_i_I clknet_4_11__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06551__I _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08051__B2 as2650.indirect_target\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11169__I _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10073__I _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07970_ _02614_ _01764_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06921_ _01803_ _01835_ _01836_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09551__A1 _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06852_ as2650.debug_psl\[2\] _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09640_ _02676_ _04318_ _04320_ _02658_ _04325_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
Xclkbuf_leaf_109_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_109_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05803_ _00796_ as2650.regs\[7\]\[3\] _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09571_ _01497_ _01614_ _01491_ _01598_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06783_ _01278_ _01703_ _01364_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_78_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08522_ _01452_ _03226_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05734_ _00662_ _00738_ _00739_ _00741_ _00746_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_91_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06117__A1 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07165__I0 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11110__A1 _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08453_ _01823_ _03164_ _03168_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05665_ as2650.insin\[1\] _00663_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_77_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__B2 _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07404_ _02062_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08384_ _03104_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_129_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05596_ as2650.PC\[2\] _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__05630__I as2650.page_reg\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09606__A2 _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07335_ net123 _02139_ _02175_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07617__A1 net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10216__A3 _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05628__B1 _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07266_ _02113_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09005_ _02919_ _03696_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_130_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06217_ _01172_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07197_ _02054_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input63_I rom_bus_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06148_ _01119_ _01105_ _01106_ _01120_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__08042__A1 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10924__A1 _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09790__A1 _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06079_ _01059_ net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_109_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09907_ _04556_ net148 _04557_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_137_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09838_ net44 as2650.irqs_latch\[1\] _04514_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_154_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09769_ _04440_ _01701_ _04451_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11800_ _00579_ clknet_leaf_25_wb_clk_i as2650.stack\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09696__I2 net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11731_ _00515_ clknet_leaf_19_wb_clk_i as2650.stack\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07856__B2 _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06636__I _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11662_ _00446_ clknet_leaf_96_wb_clk_i as2650.regs\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10613_ _05092_ _05123_ _05128_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11593_ _00377_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10544_ as2650.stack\[15\]\[2\] _05076_ _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_84_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10475_ as2650.stack\[2\]\[10\] _05033_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06831__A2 _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_7_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09781__A1 _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11027_ _01819_ _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_142_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10143__A2 _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05715__I _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07847__A1 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09300__A4 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07120_ net70 _02007_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07051_ _00722_ _01770_ _01956_ _01717_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_67_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06002_ _01001_ _01002_ _00603_ _00596_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__07377__I _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput113 net113 RAM_end_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_149_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput124 net124 RAM_start_addr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput135 net135 RAM_start_addr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput146 net146 bus_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput157 net157 bus_we_sid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09772__A1 net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput168 net168 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput179 net179 io_out[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06586__A1 _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07953_ _02711_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06904_ _01738_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07884_ _01720_ _02645_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10134__A2 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09623_ _02576_ _04306_ _04308_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06835_ _01754_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_155_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09554_ _03627_ _03636_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06766_ _01686_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07840__I _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08505_ _01689_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05717_ _00729_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_91_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07838__A1 _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06697_ _01616_ _01601_ _01624_ net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_09485_ _04170_ _04056_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_93_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05648_ _00661_ _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__06456__I _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08436_ as2650.insin\[6\] _02612_ _02463_ _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_77_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_138_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08367_ _01160_ _03088_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05579_ as2650.relative_cyc as2650.indirect_cyc as2650.cycle\[9\] as2650.is_interrupt_cycle
+ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_50_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07318_ _02130_ _02159_ _02161_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08263__A1 as2650.instruction_args_latch\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08298_ _02997_ _03024_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_134_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07249_ _02086_ net129 _02087_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10706__I _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05616__A3 _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10260_ _04166_ _04783_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _04769_ _04695_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09007__I _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09818__A2 _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07829__A1 _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11714_ _00498_ clknet_leaf_119_wb_clk_i as2650.stack\[6\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11645_ _00429_ clknet_leaf_26_wb_clk_i as2650.stack\[7\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 bus_in_serial_ports[6] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07057__A2 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput26 bus_in_timers[1] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11576_ _00360_ clknet_leaf_88_wb_clk_i as2650.stack\[3\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 io_in[4] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_13_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput48 irqs[5] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 rom_bus_in[1] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10527_ _04659_ _05065_ _05068_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10458_ _04633_ _05019_ _05025_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10389_ _04777_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_144_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08309__A2 as2650.instruction_args_latch\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06620_ _01556_ _01558_ _01563_ net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_53_1801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06740__A1 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06551_ _01263_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11182__I _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09270_ _03937_ _03954_ _03955_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06099__A3 _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07296__A2 _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06482_ _01444_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08493__A1 _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08221_ _01040_ _02950_ _02957_ _02958_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_5_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_1456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08152_ as2650.ivectors_base\[10\] _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_99_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07103_ as2650.stack\[11\]\[13\] _01993_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08424__C _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08083_ as2650.ivectors_base\[4\] _02744_ _02670_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09993__A1 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08796__A2 _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07034_ _01930_ _01940_ _01942_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06559__A1 _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_124_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_124_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_1541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07835__I _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08985_ _03673_ _03674_ _03676_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_23_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07936_ as2650.irqs_latch\[4\] _02694_ _02695_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_127_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10107__A2 _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input26_I bus_in_timers[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07867_ _02462_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_74_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09606_ _02579_ _01837_ _02471_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06818_ _01738_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06731__A1 _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07798_ _02566_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_79_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09537_ _01200_ _03677_ _04219_ _04222_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_94_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06749_ _01638_ _01671_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07503__C _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09468_ _04132_ _04149_ net218 net194 _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_94_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06495__B1 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10291__A1 _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08419_ as2650.stack\[8\]\[15\] _03137_ _03138_ as2650.stack\[9\]\[15\] _03131_ _03139_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_97_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09399_ _03977_ _03978_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11430_ _00214_ clknet_leaf_52_wb_clk_i as2650.instruction_args_latch\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08236__A1 as2650.instruction_args_latch\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06914__I _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11361_ _00157_ clknet_leaf_105_wb_clk_i wb_counter\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10312_ _01637_ _04887_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_61_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11292_ _00088_ clknet_leaf_155_wb_clk_i net277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_127_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09736__A1 _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ _01413_ _04820_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_37_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09736__B2 _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10174_ _02893_ as2650.instruction_args_latch\[14\] _02474_ _04753_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10171__I _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06722__A1 _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10282__A1 _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05828__A3 _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11628_ _00412_ clknet_leaf_20_wb_clk_i as2650.stack\[15\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10034__A1 as2650.stack\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09975__A1 _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmax_cap304 _01535_ net304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_11559_ _00343_ clknet_leaf_121_wb_clk_i as2650.stack\[10\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06789__A1 _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11437__CLK clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08950__A2 _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i clknet_4_6__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05982_ _00974_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08770_ as2650.stack\[7\]\[8\] _03466_ _03462_ as2650.stack\[6\]\[8\] _03467_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07721_ _02489_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_108_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08702__A2 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ _02384_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06713__A1 net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07390__I _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08419__C _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06603_ _01545_ clknet_1_0__leaf__01549_ net175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07583_ wb_counter\[13\] _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _04006_ _04007_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_06534_ _00874_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_87_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07269__A2 _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08466__A1 as2650.ivectors_base\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09253_ _00756_ _00791_ _01493_ _03938_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06465_ as2650.debug_psl\[6\] _01188_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_69_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08204_ _01233_ _02944_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09184_ _01023_ _00816_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06396_ _01346_ _01360_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_161_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09966__A1 _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ as2650.instruction_args_latch\[12\] _02660_ _02712_ _02884_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_117_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08066_ _02793_ _02819_ _02804_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_77_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07017_ _01783_ _01922_ _01926_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_101_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09718__A1 _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_73_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08941__A2 as2650.debug_psl\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ _01606_ net356 _03588_ _01607_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_86_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06952__A1 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_86_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07919_ _01264_ _02633_ _01472_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_output132_I net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08899_ _01855_ _03587_ _03590_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_93_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08396__I _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10930_ _04949_ _05302_ _05366_ _05367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_92_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_21_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10861_ _05275_ _05302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_168_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08457__A1 _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10792_ _05092_ _05237_ _05242_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09957__A1 net223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11413_ _00197_ clknet_leaf_71_wb_clk_i as2650.indexed_cyc\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_39_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08999__C _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11344_ net379 clknet_leaf_141_wb_clk_i wb_counter\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09709__A1 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11275_ _00071_ clknet_leaf_108_wb_clk_i net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_24_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05994__A2 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10226_ _01568_ _01614_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_101_1411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08932__A2 _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ _01503_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10088_ as2650.stack\[3\]\[5\] _04676_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10255__A1 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08999__A2 _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07120__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06250_ _01102_ _01222_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06181_ _01132_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_41_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10558__A2 _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07423__A2 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09940_ net144 _04576_ _04579_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_111_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10804__I _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07385__I _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09871_ as2650.stack\[5\]\[5\] _04534_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08822_ _03250_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_124_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08753_ _03070_ _03092_ _03094_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_05965_ _00968_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_158_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07704_ _02472_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05896_ _00589_ _00837_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08684_ as2650.stack\[15\]\[5\] _02508_ _02540_ as2650.stack\[14\]\[5\] _03204_ _03384_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__10494__A1 as2650.stack\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07635_ wb_counter\[23\] _02416_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07566_ _02363_ _02364_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_0_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09305_ _03982_ _03989_ _03990_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_53_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06517_ _01314_ _01267_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_118_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07497_ net358 _02307_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09236_ _01023_ _00792_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06448_ _01373_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_20_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07662__A2 _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08880__S _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_79_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06379_ _00778_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09167_ _03160_ _03850_ _03853_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_75_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08118_ _02788_ _01908_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08611__A1 _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09098_ _01771_ _02478_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_124_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08049_ _02803_ _02705_ _02647_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_102_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07295__I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11060_ _01946_ _05473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_134_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10011_ _02537_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06639__I _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08142__A3 _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10913_ _03362_ _05321_ _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_168_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10844_ _05147_ _05258_ _05286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_168_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_143_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ as2650.stack\[6\]\[0\] _05232_ _05233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_94_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_82_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08850__A1 as2650.stack\[8\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08850__B2 as2650.stack\[9\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05664__A1 _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11327_ net368 clknet_leaf_146_wb_clk_i web_behavior\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10624__I _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07419__B _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_152_Left_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10960__A2 _05391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11258_ _00054_ clknet_leaf_149_wb_clk_i net132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08905__A2 _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10209_ as2650.regs\[5\]\[0\] _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_158_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11189_ as2650.stack\[9\]\[3\] _05551_ _05555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10712__A2 _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05750_ _00761_ net202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_76_1483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05681_ as2650.regs\[3\]\[7\] _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_118_1782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_161_Left_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07192__I1 net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07420_ _02220_ _02248_ _02250_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_158_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08764__I _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07351_ _02078_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_70_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09094__A1 _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06302_ _01272_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06284__I _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07282_ _02080_ _02127_ _02129_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_143_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06233_ _01205_ _01195_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09021_ _03703_ _03712_ _03700_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_5_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06164_ net65 _01080_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__A2 _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05670__A4 _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09528__C _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06095_ _01062_ _01064_ _01068_ _01071_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_70_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05958__A2 as2650.instruction_args_latch\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10951__A2 _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09923_ _04562_ _01674_ _04568_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08004__I _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_127_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09854_ _01961_ _04522_ _04523_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08805_ _01480_ _01895_ _03500_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_107_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _04464_ _04466_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06997_ _01907_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08736_ _03430_ _03431_ _03432_ _03433_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05948_ _00944_ _00952_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_154_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10467__A1 as2650.stack\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08667_ _02595_ _03366_ _03367_ _03225_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05879_ _00692_ _00884_ _00885_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__07183__I1 net120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07618_ _02390_ _02405_ _02406_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_132_1757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08598_ as2650.stack\[11\]\[2\] _03289_ _03290_ as2650.stack\[10\]\[2\] _03301_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__10219__A1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07549_ _02292_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_53_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06194__I _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08832__A1 _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10560_ _01868_ _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_107_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ _03885_ _03901_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10491_ _05045_ _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09719__B _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06922__I _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09632__I0 _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07399__A1 _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08596__B1 _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__05949__A2 as2650.instruction_args_latch\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11112_ _05455_ _05502_ _05506_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11043_ _05440_ _05461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_53_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08899__A1 _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09173__C _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09699__I0 net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10458__A1 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07174__I1 net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05885__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ net219 _05266_ _05267_ _05268_ _05269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_156_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10758_ as2650.regs\[6\]\[3\] _05221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10225__A4 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10689_ _04721_ _05165_ _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_125_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11186__A2 _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08051__A2 _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06920_ as2650.stack\[12\]\[5\] _01821_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06851_ _01752_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05802_ as2650.regs\[3\]\[3\] _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09570_ _04194_ _01401_ _01768_ _01349_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_155_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06782_ _01163_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_91_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08521_ _01473_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_102_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05733_ _00745_ as2650.instruction_args_latch\[7\] _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_102_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06117__A2 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07165__I1 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_149_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_149_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08452_ as2650.ivectors_base\[1\] _03165_ _03167_ _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05664_ _00667_ _00677_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_65_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07403_ _02220_ _02234_ _02235_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05595_ as2650.cycle\[4\] as2650.indirect_target\[0\] _00598_ _00609_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09067__A1 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08383_ _01240_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09606__A3 _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07334_ _02121_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_1652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05628__A1 as2650.indirect_target\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05628__B2 as2650.page_reg\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07265_ _02112_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09004_ _03657_ _03591_ _03695_ _01462_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_162_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06216_ _01186_ _01188_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_147_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07196_ net95 net111 _02051_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06147_ net41 _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08042__A2 _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input56_I ram_bus_in[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06078_ _00841_ net353 _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09790__A2 _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09906_ _04555_ _01599_ _04558_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_6_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10137__B1 _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09837_ _01516_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_57_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09768_ _04432_ _02556_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output212_I net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08719_ _01848_ _03417_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_68_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09699_ net3 net11 net27 net19 _04383_ _04384_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__08502__B1 _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11101__A2 _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09696__I3 net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11730_ _00514_ clknet_leaf_77_wb_clk_i as2650.regs\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05821__I _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11661_ _00445_ clknet_leaf_96_wb_clk_i as2650.regs\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10612_ as2650.stack\[7\]\[7\] _05124_ _05128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08805__A1 _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11592_ _00376_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10543_ _01776_ _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07748__I _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10474_ _04649_ _05032_ _05035_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_161_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08569__B1 _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10915__A2 _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09781__A2 _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07792__A1 _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08800__C _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11026_ _05447_ _05439_ _05448_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07432__B _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06827__I _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07847__A2 _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11859_ net187 net261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_151_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09844__I0 as2650.trap vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10603__A1 _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07050_ as2650.debug_psu\[7\] _01773_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06001_ as2650.is_interrupt_cycle _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_109_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10084__I _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput114 net114 RAM_end_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_149_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput125 net125 RAM_start_addr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput136 net136 RAM_start_addr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput147 net147 bus_data_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput158 net158 bus_we_timers vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput169 net169 io_oeb[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06586__A2 _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07952_ _01250_ _01244_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_103_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__A3 _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06903_ _01819_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_103_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07883_ _00686_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_138_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08732__B1 _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ _01568_ _04307_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06834_ as2650.debug_psl\[1\] _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09553_ _04234_ _04236_ _04237_ _04238_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06765_ as2650.debug_psu\[0\] as2650.debug_psu\[1\] _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08504_ as2650.stack\[12\]\[0\] _02532_ _02535_ as2650.stack\[13\]\[0\] _03209_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05716_ _00728_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ _04025_ _04043_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06696_ net247 _01617_ _01612_ _01623_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_91_1586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ _02803_ _01337_ _03152_ _03153_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_109_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05647_ _00660_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ net209 _01438_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05578_ as2650.PC\[7\] _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_11_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07317_ net295 _02137_ _02160_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08297_ _02998_ _02637_ _03020_ _03010_ _03023_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_117_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07248_ _02084_ net160 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_95_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_46_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_46_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_131_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__A2 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _02044_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_1823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _03816_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09763__A2 _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A3 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_340 la_data_out[51] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_167_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11713_ _00497_ clknet_leaf_119_wb_clk_i as2650.stack\[6\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06501__A2 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11644_ _00428_ clknet_leaf_130_wb_clk_i as2650.stack\[7\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput16 bus_in_serial_ports[7] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_135_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09451__A1 net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11575_ _00359_ clknet_leaf_122_wb_clk_i as2650.stack\[3\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput27 bus_in_timers[2] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08083__B _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput38 io_in[5] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput49 irqs[6] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06382__I _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10526_ as2650.stack\[1\]\[13\] _05066_ _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10457_ as2650.stack\[2\]\[3\] _05021_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10388_ _02553_ _04934_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06407__I3 _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i clknet_4_5__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07427__B _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11009_ _05391_ _05398_ _05434_ _05435_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_75_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08190__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06550_ _01504_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ _01443_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06099__A4 _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08220_ _02933_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09868__I _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08151_ _02888_ _02747_ _02892_ _02898_ _02745_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_28_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07102_ _01940_ _01992_ _01994_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06256__A1 _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06292__I _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08082_ _02604_ _02834_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07033_ as2650.stack\[12\]\[12\] _01941_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06008__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05837__S _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08984_ _03675_ _03643_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07935_ as2650.irqs_latch\[5\] _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_1740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07508__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07866_ _02624_ _02629_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_88_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07851__I _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09605_ _02665_ _02470_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_input19_I bus_in_sid[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06817_ _01714_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_79_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07797_ _01183_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09536_ _03676_ _03772_ _03775_ _03613_ _04221_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_52_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06748_ _01665_ _01670_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10815__A1 _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ _04146_ _04151_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06679_ _01606_ _01598_ _01607_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_8_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09681__A1 _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06495__A1 _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08418_ _02535_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09398_ _04083_ _03927_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_97_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08349_ net209 _02575_ _03067_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_69_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10717__I _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06247__A1 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11360_ _00156_ clknet_leaf_104_wb_clk_i wb_counter\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07995__A1 _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ _04358_ _01372_ as2650.debug_psl\[5\] _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11291_ _00087_ clknet_leaf_155_wb_clk_i net266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_123_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10242_ _02913_ _02927_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_37_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10173_ _04750_ _04751_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_100_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08172__A1 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07761__I _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08078__B _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11627_ _00411_ clknet_leaf_23_wb_clk_i as2650.stack\[15\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09424__A1 _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09975__A2 _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11558_ _00342_ clknet_leaf_124_wb_clk_i as2650.stack\[10\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xmax_cap305 _00608_ net305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_53_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10509_ _04641_ _05053_ _05057_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11489_ _00273_ clknet_leaf_0_wb_clk_i as2650.stack\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06840__I _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07738__A1 as2650.stack\[0\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06410__A1 _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05981_ _00939_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07720_ _02488_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08163__A1 _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07651_ wb_counter\[27\] _02432_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06713__A2 net237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06602_ clknet_leaf_36_wb_clk_i _01548_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06287__I _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07582_ _02373_ _02375_ _02377_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_53_1643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09321_ _03969_ _03970_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_88_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06533_ _01492_ net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_158_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06477__A1 _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09252_ _00855_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06464_ _00680_ _01224_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_63_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08435__C _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08203_ _02943_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09183_ _00765_ _00888_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10537__I _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06395_ _01347_ _01348_ _01359_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06229__A1 _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08134_ as2650.indirect_target\[12\] _02680_ _02844_ _02882_ _02883_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_71_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08065_ _02816_ _02818_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_82_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07846__I _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07016_ _01924_ _01731_ _01925_ _01717_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_102_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10272__I _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_129_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06401__A1 _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08967_ _03658_ _01212_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07918_ _01702_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_86_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_1670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08898_ _03589_ _01677_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08154__A1 _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output125_I net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07849_ _02614_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_54_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06704__A2 _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10860_ _05294_ _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_151_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09519_ _03653_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09654__A1 _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10791_ as2650.stack\[6\]\[7\] _05238_ _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_72_wb_clk_i_I clknet_4_15__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09406__A1 _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11412_ _00196_ clknet_leaf_71_wb_clk_i as2650.indexed_cyc\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09957__A2 _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11343_ net375 clknet_leaf_143_wb_clk_i wb_counter\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07756__I _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11274_ _00070_ clknet_leaf_112_wb_clk_i net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_39_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10182__I _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ _01237_ _01099_ _01182_ _01169_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__09971__I _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _01411_ _01504_ _04734_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_98_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__I _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _04635_ _04675_ _04677_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__A1 _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10989_ _05347_ _05412_ _05416_ as2650.regs\[0\]\[3\] _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06459__A1 _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06835__I _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07408__B1 _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11204__A1 _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06180_ _01111_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05895__B _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06570__I _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_165_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09870_ _01820_ _04533_ _04535_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_117_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08821_ _03248_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09814__C _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ _03372_ _03427_ _03449_ _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05964_ net227 net246 _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__05914__I net200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07703_ _02466_ _02471_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_94_1754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08683_ as2650.stack\[12\]\[5\] _02532_ _02535_ as2650.stack\[13\]\[5\] _03383_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05895_ net305 _00836_ _00612_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09884__A1 _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07634_ _02407_ _02417_ _02419_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_105_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07565_ wb_counter\[9\] wb_counter\[10\] _02359_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09636__A1 _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09304_ _01024_ net220 _03987_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06516_ as2650.cycle\[10\] _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_118_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07496_ wb_reset_override_en _02305_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08165__C _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09235_ _00718_ _00826_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06447_ _01405_ _01339_ _01407_ _01409_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_118_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09166_ _01434_ _03786_ _03851_ _03852_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06378_ _00935_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_75_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08117_ _02800_ _01919_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _03737_ _03311_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08048_ _02802_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06480__I _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07509__C _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10010_ _01736_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output242_I net242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09999_ _01928_ _04609_ _04614_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08127__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08200__I _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08678__A2 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10912_ _05349_ _05297_ _05298_ _00921_ _05350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08142__A4 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09740__B _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10485__A2 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_28_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10843_ _01085_ _05284_ _05285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10774_ _05231_ _05232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09031__I _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07102__A2 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__I _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05664__A2 _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11326_ _00122_ clknet_leaf_153_wb_clk_i web_behavior\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06390__I _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11257_ _00053_ clknet_leaf_152_wb_clk_i net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08366__A1 net209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10208_ _04786_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11188_ _05445_ _05549_ _05554_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_160_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10139_ _01082_ _01573_ _03743_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_59_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08118__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08110__I as2650.instruction_args_latch\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09866__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05680_ _00693_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A1 _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ _02162_ _02186_ _02189_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06301_ _01192_ _01163_ _01213_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_143_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07281_ net291 _02095_ _02128_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08841__A2 _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09020_ _03699_ _03698_ _03705_ _03711_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06232_ _01173_ _01179_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_2_1477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold116_I wbs_dat_i[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06163_ net36 _01133_ _01135_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_14_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05909__I _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06094_ net233 net252 _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_145_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09922_ _04563_ net154 _04564_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10951__A3 _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08357__A1 _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09853_ _01901_ _01924_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10164__A1 _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10550__I _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08804_ _03197_ _03484_ _03499_ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09784_ _04465_ _01901_ _01701_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06996_ _01905_ _01906_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08109__B2 _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08735_ as2650.stack\[4\]\[7\] _03411_ _03412_ as2650.stack\[5\]\[7\] _02517_ _03433_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05947_ _00940_ _00627_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_1_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05591__A1 _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07868__B1 _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08955__I _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08666_ _01812_ _01574_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05878_ _00707_ as2650.regs\[7\]\[2\] _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07617_ net84 _02394_ _02401_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08597_ _03291_ _03295_ _03297_ _03299_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09609__A1 as2650.debug_psu\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ wb_counter\[7\] _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09704__S1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_7__f_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07096__A1 _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07479_ _02239_ wb_counter\[31\] _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09218_ _03870_ _03872_ _03903_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_63_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output192_I net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10490_ _05044_ _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_134_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09149_ _03824_ _03834_ _03835_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_60_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07399__A2 _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09632__I1 _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11111_ as2650.stack\[14\]\[6\] _05503_ _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_57_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08348__A1 _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11042_ _05438_ _05460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_53_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08899__A2 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10460__I _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09699__I1 net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold94_I wbs_dat_i[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10826_ _03218_ _05266_ _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06385__I _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09076__A2 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10757_ _05172_ _05215_ _05217_ _05220_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_153_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08823__A2 _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05637__A2 _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10630__A2 _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10688_ _05179_ _05175_ _05176_ _00710_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_153_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11309_ _00105_ clknet_leaf_105_wb_clk_i net275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09536__B1 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06850_ _01768_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05801_ _00657_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_136_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06781_ _01302_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_116_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08520_ _03224_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05732_ _00744_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_56_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06117__A3 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08511__A1 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08708__C _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08451_ _01547_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05663_ _00665_ _00675_ _00676_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_TAPCELL_ROW_19_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_11_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07402_ net275 _02225_ _02218_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08382_ _03056_ _03066_ _03100_ _03103_ _02942_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_19_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05594_ _00606_ _00593_ _00595_ _00603_ _00607_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07333_ _02115_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07078__A1 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08814__A2 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_118_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_118_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05628__A2 _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07264_ net70 _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_1528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ _03690_ _03691_ _03694_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_131_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06215_ _01187_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_144_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ _02053_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10909__B1 _05347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08578__A1 _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06146_ _01104_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06077_ net229 net248 _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_22_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09790__A3 _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07854__I _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I irqs[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09905_ _04556_ net147 _04557_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_6_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10137__A1 _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10137__B2 _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09836_ _04513_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06979_ as2650.PC\[8\] _01862_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09767_ _03141_ _03143_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_20_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08718_ _01831_ _03387_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09698_ as2650.ext_io_addr\[6\] _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_96_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08502__B2 as2650.stack\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08649_ _01475_ _02754_ _03349_ _03237_ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_output205_I net205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11660_ _00444_ clknet_leaf_78_wb_clk_i as2650.regs\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10611_ _05090_ _05123_ _05127_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11591_ _00375_ clknet_leaf_12_wb_clk_i as2650.stack\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08805__A2 _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05619__A2 _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10542_ _05078_ _05074_ _05079_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_59_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10473_ as2650.stack\[2\]\[9\] _05033_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08569__B2 _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10376__A1 _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07241__A1 _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07764__I _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i clknet_4_4__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_44_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07792__A2 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10128__A1 as2650.cycle\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11025_ as2650.stack\[0\]\[3\] _05441_ _05448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09297__A2 _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_155_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__A1 _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11858_ net298 net260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_151_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_151_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10809_ as2650.stack\[6\]\[14\] _05250_ _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11789_ _00568_ clknet_leaf_110_wb_clk_i as2650.stack\[13\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07939__I _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07480__A1 _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06000_ _00591_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput115 net115 RAM_end_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10367__A1 _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput126 net126 RAM_start_addr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput137 net137 RAM_start_addr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput148 net148 bus_data_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput159 net159 cs_port[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07951_ _02698_ _02709_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10119__A1 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06902_ _01811_ _01818_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07882_ _02643_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_120_1470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08732__B2 as2650.stack\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06833_ _01752_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09621_ _01577_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09552_ _04232_ _03773_ _03775_ _03661_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_06764_ _01684_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08503_ as2650.stack\[8\]\[0\] _02525_ _02528_ as2650.stack\[9\]\[0\] _02504_ _03208_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_56_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08438__C _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07299__A1 net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05715_ _00727_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__08496__B1 _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _04057_ _04068_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06695_ _01618_ _01622_ _01527_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_56_1696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08434_ _02595_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_93_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05646_ _00657_ _00659_ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08365_ _03074_ _03085_ _03086_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05577_ _00590_ _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_138_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07849__I _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07316_ _02074_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ _03021_ _02620_ _03022_ net207 _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_11_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07247_ wb_debug_carry _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07178_ net86 net118 _02041_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06129_ _01101_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08420__B1 _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_86_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_86_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_140_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08971__A1 _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output155_I net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_15_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_15_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08723__A1 _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09819_ _02570_ _04497_ _04498_ _03049_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_96_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07533__B _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09279__A2 _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_as2650_330 la_data_out[33] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_51_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xwrapped_as2650_341 la_data_out[52] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_96_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11712_ _00496_ clknet_leaf_89_wb_clk_i as2650.stack\[6\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06501__A3 _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11643_ _00427_ clknet_leaf_22_wb_clk_i as2650.stack\[7\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07759__I _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11574_ _00358_ clknet_leaf_123_wb_clk_i as2650.stack\[3\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10597__A1 _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 bus_in_sid[0] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09451__A2 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput28 bus_in_timers[3] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_1694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput39 io_in[6] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10185__I _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07462__A1 net285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10525_ _04655_ _05065_ _05067_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10456_ _04631_ _05019_ _05024_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_1708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09203__A2 _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08811__C _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ _04959_ _04960_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_23_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11008_ as2650.regs\[0\]\[7\] _05405_ _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06480_ _01442_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08150_ as2650.indirect_target\[13\] _02761_ _02713_ _02897_ _02718_ _02898_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_43_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07101_ as2650.stack\[11\]\[12\] _01993_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10095__I _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ _02698_ _02832_ _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06256__A2 _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07032_ _01738_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_114_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07205__A1 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11001__A2 _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _03616_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07934_ as2650.irqs_latch\[1\] _02693_ as2650.irqs_latch\[3\] _02694_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_97_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_127_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07865_ as2650.insin\[4\] _02596_ _02628_ _02600_ _02604_ _02629_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_88_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08449__B _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ _03731_ _04289_ _03721_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_155_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06816_ _01736_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07796_ _02467_ _02564_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05652__I _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06747_ _01604_ _01669_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09535_ _02467_ _04220_ _03675_ _02564_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_6_1409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11068__A2 _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_133_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_133_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09130__A1 _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09466_ _04146_ _04151_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06678_ _01043_ _01490_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10815__A2 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09681__A2 _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_4_12__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05629_ _00640_ _00642_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08417_ _02532_ _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_93_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09397_ _03902_ _03906_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_1409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08348_ _02788_ _03069_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07444__A1 net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06247__A2 _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03005_ _03008_ _02622_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10310_ _04733_ _04884_ _04885_ _04740_ _04194_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__07995__A2 _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11290_ _00086_ clknet_4_0__leaf_wb_clk_i net265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08631__C _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10241_ _04817_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_37_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_37_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10172_ _01412_ _04711_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08203__I _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_1785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06183__A1 _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11059__A2 _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__C1 _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09121__A1 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09969__I _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10806__A2 _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11626_ _00410_ clknet_leaf_20_wb_clk_i as2650.stack\[15\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09424__A2 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11557_ _00341_ clknet_leaf_125_wb_clk_i as2650.stack\[10\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ as2650.stack\[1\]\[6\] _05054_ _05057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11488_ _00272_ clknet_leaf_4_wb_clk_i as2650.stack\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10439_ _05010_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_106_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_107_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05980_ _00973_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07650_ wb_counter\[26\] _02429_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06568__I _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06601_ _01547_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_122_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07910__A2 _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07581_ net396 _02376_ _02368_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05921__A1 _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09320_ _03991_ _04004_ _04005_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09112__A1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06532_ _01491_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09251_ _03929_ _03936_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_75_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07674__A1 _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06463_ _01382_ _01417_ _01423_ _01425_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_135_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08871__B1 _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08202_ _01221_ _02597_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_146_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09182_ _03752_ _03868_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06394_ _01349_ _01358_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_16_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08133_ _01936_ _02881_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_146_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06229__A2 _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__B1 _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08064_ _02801_ _01845_ _02817_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_1763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07015_ net190 _01732_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08926__A1 _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06401__A2 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08966_ _00853_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08958__I _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input31_I bus_in_timers[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07917_ _02676_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_86_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08897_ _03588_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08154__A2 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09351__A1 net220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07848_ _02613_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_98_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_162_Right_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_3_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output118_I net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05912__A1 _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07779_ _02546_ _02547_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_71_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09103__A1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09518_ _03689_ _03652_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10790_ _05090_ _05237_ _05241_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09654__A2 _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08626__C _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10728__I _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09449_ _04133_ _04112_ _04134_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_23_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11411_ _00195_ clknet_leaf_46_wb_clk_i as2650.indirect_target\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_117_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11213__A2 _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11342_ _00138_ clknet_leaf_142_wb_clk_i wb_counter\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06941__I _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_30_wb_clk_i clknet_4_6__leaf_wb_clk_i clknet_leaf_30_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11273_ _00069_ clknet_leaf_109_wb_clk_i net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__09709__A3 _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08917__A1 _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10224_ _04795_ _04797_ _04800_ _04801_ _01747_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_63_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10724__A1 _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10155_ _04702_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10086_ as2650.stack\[3\]\[4\] _04676_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09342__A1 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10988_ _05333_ _05409_ _05418_ _05419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07408__A1 _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11609_ _00393_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06851__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08908__A1 _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08820_ as2650.stack\[3\]\[10\] _03461_ _03514_ as2650.stack\[2\]\[10\] _03515_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09581__A1 _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10191__A2 _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05963_ _00967_ net246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_124_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08751_ _03374_ _03445_ _03448_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08136__A2 _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09333__A1 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07702_ _02469_ _02470_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xclkbuf_0__01549_ _01549_ clknet_0__01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05894_ _00742_ as2650.instruction_args_latch\[2\] _00659_ _00899_ _00900_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_08682_ as2650.stack\[8\]\[5\] _02491_ _02498_ as2650.stack\[9\]\[5\] _03130_ _03382_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_120_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07633_ net87 _02410_ _02418_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07564_ wb_counter\[9\] _02359_ wb_counter\[10\] _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09636__A2 _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06515_ _01463_ _01470_ _01475_ _01247_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09303_ _03987_ _03988_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07495_ _02306_ net367 _02309_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08844__B1 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06446_ _01366_ _01408_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_118_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09234_ _03892_ _01028_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09165_ _03736_ _03386_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06377_ _01341_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08116_ _02623_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07857__I _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_39_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09096_ _03729_ _02586_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10954__A1 _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08047_ _02801_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_1570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05830__B1 _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08375__A2 as2650.instruction_args_latch\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__A1 _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09998_ as2650.stack\[4\]\[11\] _04610_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08949_ _00833_ _01226_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_48_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_51_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10911_ _04929_ _04930_ _05349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_28_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07541__B _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10842_ _01807_ _04699_ _05283_ _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_55_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10773_ _05228_ _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_149_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__B net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11198__A1 _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07767__I _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11325_ _00121_ clknet_leaf_151_wb_clk_i wb_debug_carry vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11256_ _00052_ clknet_leaf_151_wb_clk_i net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_142_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09563__A1 _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _04700_ _04722_ _04770_ _04571_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_11187_ as2650.stack\[9\]\[2\] _05551_ _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10138_ _04716_ _04715_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_66_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07435__C _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10142__B _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10069_ _04663_ _04656_ _04664_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07007__I _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09618__A2 _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08826__B1 _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06300_ _01248_ _01271_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_75_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07280_ _02074_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06231_ _01203_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_142_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06162_ _01134_ _01133_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold109_I wbs_dat_i[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06093_ _01070_ net252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_125_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09921_ _04562_ _01664_ _04567_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09852_ _02534_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08803_ _01445_ _03486_ _03498_ _03312_ _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08301__I _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09783_ _01682_ _03514_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06995_ as2650.PC\[8\] _01890_ _01861_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08109__A2 _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08734_ as2650.stack\[7\]\[7\] _03428_ _03429_ as2650.stack\[6\]\[7\] _03432_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05946_ _00940_ _00627_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05591__A2 _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11113__A1 as2650.stack\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05877_ as2650.regs\[3\]\[2\] _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08665_ _01816_ _03351_ _03362_ _03059_ _03365_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__07868__B2 _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07616_ wb_counter\[20\] _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_163_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_113_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08596_ as2650.stack\[4\]\[2\] _03292_ _03293_ as2650.stack\[5\]\[2\] _03298_ _03299_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09609__A2 _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_93_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07547_ wb_counter\[4\] wb_counter\[5\] wb_counter\[6\] _02336_ _02349_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_64_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07478_ as2650.wb_hidden_rom_enable _02271_ _02245_ net112 _02272_ _02298_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_107_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09217_ _00767_ net189 _03873_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_88_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06429_ _01389_ _01391_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06491__I _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ _03640_ _03615_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output185_I net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08596__A2 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09793__A1 _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ _03768_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_124_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _05453_ _05502_ _05505_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i clknet_4_3__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_57_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11041_ _01882_ _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_53_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07020__A2 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07159__I0 net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09699__I2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06126__A4 _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10825_ _05256_ _05267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10756_ as2650.regs\[6\]\[2\] _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_153_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10687_ _05011_ _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_35_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05893__I0 _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11308_ _00104_ clknet_leaf_105_wb_clk_i net274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11239_ _00035_ clknet_leaf_7_wb_clk_i as2650.stack\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07011__A2 _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05800_ _00809_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_78_1569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06780_ _01700_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_165_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05731_ _00743_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_136_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10303__C1 _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05662_ _00668_ net51 _00670_ _00672_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XTAP_TAPCELL_ROW_19_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08450_ _01804_ _03164_ _03166_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06576__I _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06522__A1 _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07401_ _02211_ wb_counter\[18\] _02233_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08381_ _03102_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_50_1411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05593_ as2650.indirect_target\[1\] _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_15_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ _02162_ _02172_ _02173_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09887__I _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _02080_ _02110_ _02111_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06525__B _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06214_ _00706_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09002_ _03692_ _03693_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08027__A1 as2650.indirect_target\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07194_ net93 net110 _02051_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07200__I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06145_ _01104_ net53 _01105_ _01106_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__08578__A2 _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09775__A1 _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06076_ _01057_ net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07250__A2 _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09527__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09904_ _03174_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_6_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10137__A2 _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09835_ _03105_ _04512_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08966__I _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ _02472_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06978_ as2650.PC\[9\] _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07870__I _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08717_ _03408_ _03415_ _02548_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05929_ _00907_ _00930_ _00931_ _00933_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_09697_ as2650.ext_io_addr\[7\] _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_69_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08502__A2 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08648_ _01475_ _01816_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08579_ _03280_ _03281_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ as2650.stack\[7\]\[6\] _05124_ _05127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_46_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11590_ _00374_ clknet_leaf_12_wb_clk_i as2650.stack\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10541_ as2650.stack\[15\]\[1\] _05076_ _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08018__A1 _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10472_ _04645_ _05032_ _05034_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_59_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09746__B _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09037__I _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11024_ _01800_ _05447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_21_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07780__I _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10420__B _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ net300 net259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_151_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10808_ _05108_ _05249_ _05252_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11788_ _00567_ clknet_leaf_132_wb_clk_i as2650.stack\[13\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10739_ as2650.stack\[8\]\[12\] _05209_ _05210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09757__A1 _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_149_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput116 net116 RAM_end_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput127 net127 RAM_start_addr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput138 net138 WEb_ram vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_161_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput149 net149 bus_data_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_142_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09509__A1 net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07950_ _00611_ _02635_ _02707_ _02708_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_103_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10119__A2 _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06901_ _01813_ _01741_ _01817_ _01798_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_07881_ _02642_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08732__A2 _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09620_ _01092_ _03720_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06832_ _01751_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09551_ _01703_ _03635_ _03632_ _01231_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_116_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06763_ _01682_ _01683_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08502_ as2650.stack\[11\]\[0\] _03200_ _02511_ as2650.stack\[10\]\[0\] _03207_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_37_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05714_ _00724_ as2650.regs\[4\]\[7\] _00726_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_06694_ _01544_ _01621_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09482_ _04070_ _04078_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08433_ _03151_ _01578_ _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05645_ _00658_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_65_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05576_ _00589_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08364_ _02625_ _03072_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_138_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ _02155_ wb_counter\[7\] _02158_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08295_ _03001_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07246_ _02080_ _02093_ _02096_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _02043_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input61_I rom_bus_in[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06128_ _01100_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06059_ _00745_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output148_I net148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09818_ _01931_ _02628_ _02589_ _03818_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_91_wb_clk_i_I clknet_4_10__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06734__A1 net244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_55_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_55_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10530__A2 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08629__C _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09749_ _01700_ _04432_ _02557_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_97_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_320 la_data_out[41] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_331 la_data_out[34] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_97_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_342 la_data_out[53] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__10294__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11711_ _00495_ clknet_leaf_124_wb_clk_i as2650.stack\[6\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11642_ _00426_ clknet_leaf_22_wb_clk_i as2650.stack\[7\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11573_ _00357_ clknet_leaf_129_wb_clk_i as2650.stack\[3\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput18 bus_in_sid[1] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 bus_in_timers[4] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10524_ as2650.stack\[1\]\[12\] _05066_ _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10455_ as2650.stack\[2\]\[2\] _05021_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07214__A2 _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10386_ _04216_ _04726_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_144_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09990__I _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11007_ _05397_ _05433_ _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08478__A1 _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09675__B1 _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10285__A1 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05700__A2 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10037__A1 as2650.stack\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_136_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07100_ _01974_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08080_ as2650.instruction_args_latch\[8\] _01702_ _02656_ as2650.indirect_target\[8\]
+ _02653_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_71_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06256__A3 _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07031_ _01939_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_141_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08402__A1 _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_90_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ _03670_ _03671_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_80_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07933_ as2650.irqs_latch\[2\] _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_122_1599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_127_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07864_ _02627_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_39_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09603_ _01664_ _04288_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06815_ _01718_ _01726_ _01735_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_07795_ _02563_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_30_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09534_ _03613_ _03615_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08469__A1 _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06746_ _01666_ _01667_ _01668_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_155_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10995__B _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09130__A2 _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09465_ _04149_ _04150_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_91_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06677_ _01605_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08416_ as2650.stack\[11\]\[15\] _02539_ _02542_ as2650.stack\[10\]\[15\] _03136_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_168_1703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05628_ as2650.indirect_target\[15\] _00635_ _00641_ as2650.page_reg\[2\] _00642_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09396_ _03972_ _03980_ _04008_ _04080_ _04081_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_148_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_97_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08347_ net211 _01438_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_102_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_102_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08278_ _03007_ as2650.instruction_args_latch\[8\] _01256_ _03008_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07444__A2 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07229_ _02079_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_61_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10240_ _04817_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_131_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10171_ _04719_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08172__A3 _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__A2 _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09657__B1 _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09657__C2 _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07683__A2 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11625_ _00409_ clknet_leaf_33_wb_clk_i as2650.stack\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07435__A2 _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11556_ _00340_ clknet_leaf_127_wb_clk_i as2650.stack\[10\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__A1 _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10507_ _04639_ _05053_ _05056_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11487_ _00271_ clknet_leaf_2_wb_clk_i as2650.stack\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10438_ _05006_ _05008_ _05009_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_20_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10369_ _04795_ _04941_ _04942_ _04801_ _01823_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__10742__A2 _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08699__A1 _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06849__I _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06600_ _01546_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_125_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_122_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07580_ _02322_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05921__A2 _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10258__A1 _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09112__A2 _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06531_ _01490_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07901__C _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_0_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_0_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_1667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09250_ _03934_ _03935_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_118_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06462_ _01424_ _01165_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08201_ _01749_ _01223_ _02941_ _01295_ _02942_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_44_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06393_ _01353_ _01357_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09181_ _01570_ _03049_ _03800_ _03850_ _03867_ _03765_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_8_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08132_ _02789_ _01908_ _02880_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10430__A1 _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08063_ _02795_ _02798_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_109_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07014_ _01923_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_77_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08304__I as2650.instruction_args_latch\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_1639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08965_ _03582_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_32_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07916_ _02675_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_86_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08896_ _03585_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input24_I bus_in_sid[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08154__A3 _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09351__A2 _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ _01110_ _01112_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_135_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_1694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07362__A1 net126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07778_ _01681_ _02515_ as2650.debug_psu\[3\] _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09517_ _03689_ _03685_ _03687_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06729_ net250 _01078_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09448_ net194 _01025_ _04132_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_26_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _04051_ _04052_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_23_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11410_ _00194_ clknet_leaf_48_wb_clk_i as2650.indirect_target\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_23_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08614__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11341_ _00137_ clknet_leaf_147_wb_clk_i wb_counter\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10421__B2 _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10972__A2 _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11272_ _00068_ clknet_leaf_109_wb_clk_i net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_123_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10223_ _04739_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_70_wb_clk_i clknet_4_13__leaf_wb_clk_i clknet_leaf_70_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_30_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10154_ _04732_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_98_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06669__I _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10085_ _04669_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10987_ _03813_ as2650.regs\[4\]\[3\] _02669_ _05418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_112_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05667__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11608_ _00392_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__A2 net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_122_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _00323_ clknet_leaf_137_wb_clk_i as2650.stack\[4\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_111_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10715__A2 _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ _03228_ _03446_ _03447_ _03064_ _03230_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05962_ _00651_ _00966_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_124_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07701_ _01276_ _01193_ _01216_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08681_ as2650.stack\[11\]\[5\] _03200_ _01967_ as2650.stack\[10\]\[5\] _03381_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_75_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05893_ _00886_ _00889_ net197 _00898_ net345 _00703_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_139_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ _02384_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_1729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_1778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07563_ _02358_ _02360_ _02362_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_66_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09302_ _01024_ _01016_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06514_ _01474_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07494_ _02062_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07203__I _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05658__A1 net225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_1831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09233_ _03896_ _03917_ _03918_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06445_ _01405_ _01374_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_118_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_79_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09164_ _01569_ _02478_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06376_ _01281_ _01339_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_44_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09558__C _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08115_ _02624_ _02865_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10403__A1 _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10564__I _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07359__B _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09095_ _03693_ _03783_ _03784_ _03764_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_128_1561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08034__I _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08046_ _02800_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i clknet_4_2__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09572__A2 _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _01913_ _04609_ _04613_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _03611_ _03612_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09324__A2 _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output130_I net130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _03568_ _03569_ _03570_ _03571_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07335__A1 net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10910_ _05295_ _05334_ _05348_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10841_ _05141_ _05164_ _05283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09088__A1 _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10772_ _05229_ _05230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08835__A1 _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09468__C net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08063__A2 _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10407__C _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ _00120_ clknet_leaf_151_wb_clk_i wb_debug_cc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11255_ _00051_ clknet_leaf_152_wb_clk_i net129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07783__I _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10206_ _04780_ _04784_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_66_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11186_ _05443_ _05549_ _05553_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08771__B1 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10137_ _01182_ _01169_ _01425_ _01442_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_1729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10068_ as2650.stack\[10\]\[15\] _04657_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_130_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06230_ _01103_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11189__A2 _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06161_ net57 _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_143_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06065__A1 _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06092_ _01036_ _01069_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_48_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09920_ _04563_ net153 _04564_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_70_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07693__I _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09851_ _04521_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08802_ _03491_ _03497_ _02551_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09782_ _04451_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06994_ as2650.PC\[10\] _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08733_ as2650.stack\[0\]\[7\] _03411_ _03412_ as2650.stack\[1\]\[7\] _02502_ _03431_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05945_ _00944_ as2650.instruction_args_latch\[8\] _00949_ _00950_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_119_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08664_ _03284_ _03364_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05876_ _00858_ _00880_ _00882_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_55_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07615_ _02403_ _02399_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__05879__A1 _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08595_ _02518_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_76_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07546_ _02341_ _02347_ _02348_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05894__A4 _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07477_ _02238_ _02296_ _02297_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09216_ _03885_ _03901_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_63_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06428_ _01390_ _01359_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ _03831_ _03832_ _03833_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06359_ _01323_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09242__A1 _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09078_ _01748_ _01703_ _02581_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_60_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output178_I net178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08029_ _02611_ _02783_ _02784_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_57_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11040_ _05457_ _05450_ _05458_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07556__A1 _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_53_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07159__I1 net127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11104__A2 _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10469__I _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_93_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10824_ _05265_ _05266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_138_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10755_ _05171_ _05215_ _05217_ _05219_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_153_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_153_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06295__A1 _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10686_ _05178_ _05175_ _05176_ _00759_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_82_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05893__I1 _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11040__A1 _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11307_ _00103_ clknet_leaf_106_wb_clk_i net273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07219__S _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09536__A2 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11238_ _00034_ clknet_leaf_7_wb_clk_i as2650.stack\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11169_ _05523_ _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07018__I _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05730_ _00742_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_117_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10303__B1 _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05661_ _00669_ _00671_ _00673_ _00674_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_19_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_4_5__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07400_ _02212_ _02231_ _02232_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_19_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08380_ _03101_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05592_ as2650.PC\[1\] _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_89_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07331_ net297 _02166_ _02160_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold121_I wbs_dat_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07262_ net288 _02095_ _02075_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09001_ _03582_ _03591_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06213_ _01185_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_144_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07193_ _02052_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10909__A2 _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11031__A1 _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06144_ _00664_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09775__A2 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__C _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06075_ _00883_ _00905_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_83_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09903_ as2650.cycle\[1\] _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_127_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_127_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09834_ _02570_ _04508_ _04511_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09765_ _04428_ _04448_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06977_ _01351_ _01753_ _01888_ _01840_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_38_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08468__B _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _03409_ _03410_ _03413_ _03414_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05928_ _00932_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06767__I _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09696_ net2 net26 net10 net18 as2650.ext_io_addr\[6\] _01518_ _04382_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_96_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08647_ _01816_ _03347_ _03194_ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10845__A1 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05859_ as2650.regs\[2\]\[1\] _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_136_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09838__I0 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08578_ _03237_ _01765_ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07529_ _02332_ _02333_ net433 _02236_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_46_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07598__I _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10540_ _01759_ _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_68_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08018__A2 _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10471_ as2650.stack\[2\]\[8\] _05033_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_157_Right_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07777__A1 _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05846__I _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07529__A1 _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10128__A3 _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11023_ _05445_ _05439_ _05446_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_142_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09053__I _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10199__I _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10836__A1 _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11856_ net184 net258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08892__I _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10807_ as2650.stack\[6\]\[13\] _05250_ _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11787_ _00566_ clknet_leaf_150_wb_clk_i as2650.stack\[13\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_126_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07465__B1 _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10738_ _05190_ _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_137_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10669_ _01240_ _05168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_152_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09757__A2 _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput106 net106 RAM_end_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput117 net117 RAM_end_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_45_1547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput128 net128 RAM_start_addr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput139 net139 boot_rom_en vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_142_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05756__I _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A1 _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09509__A2 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _01725_ _01816_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07880_ _01435_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06831_ _01749_ _01750_ _01700_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_159_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09550_ _03823_ _03664_ _04235_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06762_ as2650.debug_psu\[3\] _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08501_ _03201_ _03202_ _03203_ _03205_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_37_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10827__A1 net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05713_ _00691_ _00725_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09481_ _04008_ _04080_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_133_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06693_ _01620_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09693__A1 _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08496__A2 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08432_ _01424_ _01282_ _01198_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_153_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05644_ as2650.indexed_cyc\[1\] as2650.indexed_cyc\[0\] _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08508__S _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08735__C _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08363_ _03076_ _03082_ _03084_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_05575_ _00588_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_138_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07314_ _02116_ _02156_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_18_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07456__B1 _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08294_ _01265_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07211__I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ net266 _02095_ _02075_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_1648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07176_ net85 net117 _02041_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09566__C _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06127_ _01099_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_14_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07367__B _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08420__A2 _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input54_I ram_bus_in[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06058_ as2650.instruction_args_latch\[0\] _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06982__A2 _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08184__A1 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07881__I _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09920__A2 net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09817_ _01931_ _02480_ _04496_ _02483_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_96_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09748_ _03735_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_154_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output210_I net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10818__A1 _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_310 io_oeb[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_69_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09679_ _03783_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_119_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_321 la_data_out[42] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09684__A1 _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11710_ _00494_ clknet_leaf_22_wb_clk_i as2650.stack\[6\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xwrapped_as2650_332 la_data_out[35] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xclkbuf_leaf_95_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_95_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_343 la_data_out[54] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_55_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_24_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_24_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11641_ _00425_ clknet_leaf_40_wb_clk_i as2650.stack\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08217__I _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11572_ _00356_ clknet_leaf_127_wb_clk_i as2650.stack\[3\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 bus_in_sid[2] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07998__B2 _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10523_ _05047_ _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_1547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10454_ _04629_ _05019_ _05023_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06960__I _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10385_ _04956_ _04957_ _04958_ _04831_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__05576__I _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06422__A1 _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06973__A2 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11006_ _05011_ _05399_ _05432_ _05433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09911__A2 net150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06725__A2 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09675__A1 _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08478__A2 _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09675__B2 _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08836__B _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09978__A2 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07031__I _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_133_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08571__B _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ _01933_ _01938_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_148_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06870__I as2650.PC\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08402__A2 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08981_ _03668_ _03669_ _03672_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07932_ as2650.irqs_latch\[6\] _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08166__A1 as2650.ivectors_base\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07863_ _02626_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09602_ _01361_ _04287_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06814_ _01558_ _01731_ _01733_ _01734_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_88_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_88_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07794_ _01528_ _01151_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07206__I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09533_ _03833_ _03831_ _03832_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_30_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06745_ _01666_ _01419_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_84_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09464_ _00727_ _00722_ _04132_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_94_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06676_ _01043_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_159_Left_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08415_ _03129_ _03132_ _03133_ _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_87_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05627_ _00628_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_43_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09395_ _04006_ _04007_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_43_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08346_ net212 _02991_ _03067_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_62_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08277_ _03006_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__I _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07228_ _02078_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_127_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_142_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_142_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07159_ net77 net127 _02030_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_168_Left_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10170_ _04239_ _04729_ _04745_ _04748_ _04711_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XTAP_TAPCELL_ROW_37_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output160_I net160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_max_cap304_I _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09657__A1 _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11861__I net299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06955__I _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09409__B2 _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11624_ _00408_ clknet_leaf_33_wb_clk_i as2650.stack\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08093__B1 _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11555_ _00339_ clknet_leaf_125_wb_clk_i as2650.stack\[10\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10506_ as2650.stack\[1\]\[5\] _05054_ _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06643__A1 _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11486_ _00270_ clknet_leaf_49_wb_clk_i as2650.irqs_latch\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10437_ _04365_ _04830_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_150_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10368_ _04798_ _04737_ _01387_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10299_ _04778_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08148__A1 _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08410__I _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08699__A2 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09648__A1 _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ _01489_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_92_1684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06461_ _01277_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_8_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08871__A2 _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08200_ _01525_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_5_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_1370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06882__A1 _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09180_ _03767_ _03863_ _03866_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06392_ _01354_ _01355_ _01356_ _00853_ _01185_ _01187_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08131_ _02789_ _02877_ _02879_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08623__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__A1 _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08062_ _02787_ _01864_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_TAPCELL_ROW_12_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i clknet_4_1__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_70_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07013_ _01683_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_129_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_129_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08964_ _01462_ _03592_ _03655_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__08139__A1 _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07915_ _00678_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08895_ _03586_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08934__I0 _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07846_ _01102_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08154__A4 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05880__S _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I bus_in_sid[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _01687_ _02545_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09639__A1 _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09639__B2 _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06728_ _01649_ _01652_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09516_ _03653_ _03688_ _04200_ _04201_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_116_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09447_ _00721_ _01025_ _04132_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06659_ _01583_ _00178_ _01591_ _00180_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_82_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08862__A2 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _04051_ _04052_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_81_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_23_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08329_ _03048_ _03050_ _03051_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09811__A1 _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09811__B2 _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11340_ _00136_ clknet_leaf_146_wb_clk_i wb_counter\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11271_ _00067_ clknet_leaf_109_wb_clk_i net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_105_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08378__A1 _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10222_ _04798_ _04799_ _01415_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11856__I net184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07050__A1 as2650.debug_psu\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _01082_ _01572_ _04715_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__10760__I _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05600__A2 _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10084_ _04667_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10488__A2 _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_139_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10986_ _05408_ _05415_ _05417_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09061__I _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07105__A2 _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10000__I _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11607_ _00391_ clknet_leaf_13_wb_clk_i as2650.stack\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07408__A3 _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09802__A1 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11538_ _00322_ clknet_leaf_137_wb_clk_i as2650.stack\[4\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_169_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11469_ _00253_ clknet_leaf_59_wb_clk_i as2650.debug_psl\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_169_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08369__A1 _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09566__B1 _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10176__A1 _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05764__I _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I bus_in_serial_ports[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05961_ _00656_ _00956_ _00965_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_124_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07700_ _02468_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_79_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08680_ _03376_ _03377_ _03378_ _03379_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_1735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09680__B _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05892_ _00897_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07344__A2 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07631_ wb_counter\[23\] _02416_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_45_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06595__I _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07562_ net404 _02361_ _02351_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_1470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09097__A2 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ _03983_ _03984_ _03986_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_66_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06528__C _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06513_ _01473_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_1454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07493_ net366 _02307_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__A2 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _03897_ _03898_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_57_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05658__A2 net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06444_ _01400_ _01406_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06855__A1 _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_20_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09163_ _03849_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06375_ _01339_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05939__I _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08114_ as2650.ivectors_base\[6\] _02852_ _02864_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06607__A1 _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09094_ _03592_ _03783_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08045_ _01147_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_114_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05830__A2 as2650.instruction_args_latch\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09996_ as2650.stack\[4\]\[10\] _04610_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08780__A1 _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05594__A1 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ _03627_ _03636_ _03638_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_58_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08878_ as2650.stack\[15\]\[12\] _03466_ _03246_ as2650.stack\[14\]\[12\] _03520_
+ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_51_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07335__A2 _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output123_I net123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07829_ _01100_ _01286_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10840_ _05263_ _05277_ _05281_ _05282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_36_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10771_ _05228_ _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08426__S _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11323_ _00119_ clknet_leaf_141_wb_clk_i wb_feedback_delay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06074__A2 _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11254_ _00050_ clknet_leaf_151_wb_clk_i net122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09012__A2 _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10205_ _04167_ _04783_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07023__A1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11185_ as2650.stack\[9\]\[1\] _05551_ _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08771__A1 as2650.stack\[4\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ _01208_ _04185_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08771__B2 as2650.stack\[5\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10067_ _01958_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10330__A1 _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__A2 _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _05143_ _05283_ _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_128_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06837__A1 _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10633__A2 _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06301__A3 _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06160_ _01132_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_113_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10397__B2 _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_74_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07262__A1 net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06091_ _00810_ _00934_ _00784_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09003__A2 _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09850_ net49 as2650.irqs_latch\[7\] _01516_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_4_12__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08762__A1 _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08801_ _03492_ _03493_ _03494_ _03496_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06993_ _01369_ _01753_ _01903_ _01734_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09781_ _01902_ _01288_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05944_ _00740_ _00622_ _00948_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08732_ as2650.stack\[3\]\[7\] _03428_ _03429_ as2650.stack\[2\]\[7\] _03430_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_94_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_1652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08514__A1 _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09711__B1 _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08663_ _01813_ _03363_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05875_ _00859_ _00881_ _00879_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__10321__A1 _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07614_ wb_counter\[19\] _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08594_ as2650.stack\[7\]\[2\] _03289_ _03296_ as2650.stack\[6\]\[2\] _03297_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_132_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07545_ net390 _02344_ _02330_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08754__B _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07476_ net289 _02079_ _02293_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06427_ _01348_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_29_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09215_ _03890_ _03900_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06274__B _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _03616_ _03643_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_133_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06358_ _01317_ _01322_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08045__I _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10388__A1 _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09242__A2 _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07789__C1 _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07253__A1 _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09077_ _03701_ _03766_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06289_ _01260_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09793__A3 _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_49_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08028_ as2650.ivectors_base\[1\] _02610_ _01548_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_57_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09979_ _01801_ _04596_ _04602_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10312__A1 _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10823_ _01749_ _01728_ _02476_ _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_116_wb_clk_i_I clknet_4_9__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_1661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10754_ as2650.regs\[6\]\[1\] _05219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_82_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10685_ _04986_ _05178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05893__I2 net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_166_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11306_ _00102_ clknet_leaf_139_wb_clk_i net272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11237_ _00033_ clknet_leaf_157_wb_clk_i as2650.stack\[11\]\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08744__A1 _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11168_ _05521_ _05541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_8_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10119_ _01606_ _04697_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11099_ as2650.stack\[14\]\[1\] _05497_ _05499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_106_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_155_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05660_ net39 _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_102_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05591_ _00602_ _00594_ _00596_ _00603_ _00604_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_19_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07330_ _02155_ wb_counter\[9\] _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07261_ _02082_ _02107_ _02109_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08680__B1 _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09000_ _03592_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_166_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06212_ _00736_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_115_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold114_I wbs_adr_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07192_ net92 net109 _02051_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06143_ _01103_ _01115_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06074_ net228 _01055_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_93_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10790__A1 _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09902_ _04554_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07209__I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06113__I _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09833_ _01306_ _02589_ _04404_ _04510_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__10542__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09764_ _04446_ _04447_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06976_ _01887_ _01756_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08715_ as2650.stack\[15\]\[6\] _01687_ _01963_ as2650.stack\[14\]\[6\] _02516_ _03414_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_154_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05927_ _00925_ _00929_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11098__A2 _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09695_ _04371_ _04376_ _04379_ _04380_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_59_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08646_ _03191_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05858_ _00865_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07710__A2 _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08577_ _03192_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05789_ net201 _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_77_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07528_ net97 _02320_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_46_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07474__A1 net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07459_ _02277_ _02281_ _02283_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08671__B1 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10238__C _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output190_I net190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10470_ _05020_ _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output288_I net288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07226__A1 wb_feedback_delay vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11022__A2 _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09129_ _03816_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_103_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11022_ as2650.stack\[0\]\[2\] _05441_ _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06023__I _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06958__I _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05960__A1 _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10836__A2 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_155_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A2 _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11855_ net183 net257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_hold92_I wbs_dat_i[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10806_ _05104_ _05249_ _05251_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11786_ _00565_ clknet_leaf_133_wb_clk_i as2650.stack\[13\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10737_ _05188_ _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10668_ _05166_ _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_148_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10599_ _05078_ _05116_ _05120_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput107 net107 RAM_end_addr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_45_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput118 net118 RAM_end_addr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput129 net129 RAM_start_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_131_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09953__B _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__A3 net215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06830_ _01696_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06868__I _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07940__A2 _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ _01681_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05951__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08500_ as2650.stack\[4\]\[0\] _02525_ _02528_ as2650.stack\[5\]\[0\] _03204_ _03205_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_56_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05712_ as2650.regs\[0\]\[7\] _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_144_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06692_ _01044_ _01353_ _01619_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09480_ _03972_ _03980_ _04165_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_8_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05643_ as2650.cycle\[9\] _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08431_ _03128_ _03148_ _03150_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08362_ _02725_ _03083_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05574_ as2650.cycle\[9\] _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07313_ net182 _02141_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_138_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08293_ as2650.instruction_args_latch\[11\] _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_15_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08653__B1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07244_ _02094_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_73_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07208__A1 _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07175_ _02042_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06126_ _01098_ _00969_ _00998_ _01075_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_41_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10763__A1 _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06057_ net234 _01038_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_121_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout301 net302 net301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input47_I irqs[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08479__B _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_35_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09816_ _01804_ _02485_ _04495_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_1701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_35_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07931__A2 _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _02560_ _04429_ _04430_ _01453_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_119_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06959_ as2650.debug_psu\[0\] _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10818__A2 _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09678_ _04210_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_TAPCELL_ROW_48_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_311 io_oeb[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_48_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_as2650_322 la_data_out[43] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_333 la_data_out[36] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA_output203_I net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08629_ as2650.stack\[8\]\[3\] _03292_ _03293_ as2650.stack\[9\]\[3\] _03294_ _03331_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_96_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_344 la_data_out[55] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_84_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11640_ _00424_ clknet_leaf_40_wb_clk_i as2650.stack\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11571_ _00355_ clknet_leaf_124_wb_clk_i as2650.stack\[3\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_64_wb_clk_i clknet_4_12__leaf_wb_clk_i clknet_leaf_64_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_52_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10522_ _05045_ _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_135_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11859__I net187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10453_ as2650.stack\[2\]\[1\] _05021_ _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08233__I _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10384_ _04388_ _04764_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_60_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_144_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10506__A1 as2650.stack\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11005_ _02201_ as2650.regs\[4\]\[7\] _02669_ _05432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06688__I _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06186__A1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09064__I _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10431__C _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10809__A2 _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09675__A2 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06489__A2 _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10159__B _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11769_ _00548_ clknet_leaf_3_wb_clk_i as2650.stack\[14\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10993__A1 _05359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__I _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08938__A1 _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08980_ _03670_ _03671_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__I _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07931_ as2650.indirect_target\[1\] _02573_ _02690_ _02630_ _02691_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_23_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09363__A1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07862_ _02625_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_127_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_127_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09601_ _03732_ _03745_ _03663_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06813_ _01711_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_88_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07793_ _01263_ _01244_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_TAPCELL_ROW_88_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09115__A1 _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09532_ _03833_ _04217_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_116_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06744_ _00764_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_116_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08746__C _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06675_ _01543_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09463_ _04147_ _04148_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10848__I _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08414_ as2650.stack\[4\]\[15\] _02527_ _02530_ as2650.stack\[5\]\[15\] _03117_ _03134_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05626_ _00638_ _00639_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09394_ _04070_ _04078_ _04079_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_19_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07222__I _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07429__A1 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08345_ _01439_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08626__B1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08276_ _01307_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07227_ _02077_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_131_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_1570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _02032_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10736__A1 _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06109_ _01081_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_112_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07089_ _01972_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_100_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09593__B _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07892__I _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output153_I net153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_111_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_111_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11161__A1 _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09657__A2 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06340__A1 _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11623_ _00407_ clknet_leaf_23_wb_clk_i as2650.stack\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11216__A2 _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06971__I _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11554_ _00338_ clknet_leaf_127_wb_clk_i as2650.stack\[10\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__C _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10493__I _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10505_ _04635_ _05053_ _05055_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11485_ _00269_ clknet_leaf_49_wb_clk_i as2650.irqs_latch\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_1519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10436_ _04763_ _05007_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10367_ _04282_ _04796_ _04883_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_143_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10298_ _03528_ _04775_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08148__A2 _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06159__A1 _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09648__A2 _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10668__I _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08320__A2 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06460_ _01418_ _01340_ _01398_ _01420_ _01422_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_29_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_1394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06391_ net195 _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_50_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08130_ _02857_ _02878_ _02855_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_141_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10966__A1 _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08061_ _02814_ _02661_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_12_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_12_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07012_ _01916_ _01741_ _01921_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08802__S _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09584__A1 as2650.debug_psl\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_129_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08963_ _03582_ _03591_ _03654_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_166_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07914_ _02673_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_32_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08894_ _03585_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07198__I0 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06121__I _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07845_ _02610_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_155_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _01681_ as2650.debug_psu\[3\] _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_135_1737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09515_ _03686_ _03650_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06727_ _01544_ _01651_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10578__I _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08847__B1 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08048__I _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09446_ _04110_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06658_ _01592_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05609_ _00615_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09377_ _03997_ _03999_ _04062_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_06589_ _01537_ net164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_23_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08328_ _01087_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08075__A1 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07822__A1 _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ _02974_ _02990_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_144_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11202__I _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11270_ _00066_ clknet_leaf_109_wb_clk_i net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_127_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _04703_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10152_ _04730_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput290 net290 wbs_dat_o[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09327__A1 _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10083_ _04633_ _04668_ _04674_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07189__I0 net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07127__I _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06031__I _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07571__B _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10985_ _05330_ _05412_ _05416_ as2650.regs\[0\]\[2\] _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_70_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_27_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06313__A1 _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11606_ _00390_ clknet_leaf_13_wb_clk_i as2650.stack\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09802__A2 _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07813__A1 _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11537_ _00321_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11468_ _00252_ clknet_leaf_60_wb_clk_i as2650.debug_psl\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09566__A1 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10419_ _03744_ _04796_ _04883_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_46_1473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11399_ _00183_ clknet_leaf_49_wb_clk_i as2650.indirect_target\[3\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__10176__A2 _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08421__I _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05960_ _00961_ _00964_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_124_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05891_ _00896_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_85_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10333__C1 _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07630_ _02415_ _02412_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06552__A1 _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07561_ _02322_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08829__B1 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09300_ _03985_ _03931_ _00898_ _00875_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_66_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06512_ _01278_ _01323_ _01472_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_158_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07492_ _02146_ _02239_ _02007_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_0_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09231_ _03897_ _03898_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_88_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06443_ _01405_ _01358_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06374_ _01338_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_12_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09162_ _03764_ _03848_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10347__B _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08113_ _02837_ _02860_ _02862_ _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_126_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09093_ _03782_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _02795_ _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09006__B1 _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09557__A1 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09995_ _01899_ _04609_ _04612_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08946_ _03637_ _03626_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06791__A1 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08877_ as2650.stack\[12\]\[12\] _02492_ _02499_ as2650.stack\[13\]\[12\] _03570_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_4_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07828_ _02595_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_4_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output116_I net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ _02496_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_106_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10770_ _05016_ _04622_ _04523_ _05228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08296__B2 net207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09429_ _04114_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11322_ _00118_ clknet_leaf_140_wb_clk_i net290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_127_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11253_ _00049_ clknet_leaf_54_wb_clk_i as2650.relative_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_107_1658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _04782_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_164_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08241__I _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11184_ _05436_ _05549_ _05552_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11519__D _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10135_ _04697_ _04708_ _04709_ _04713_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__08771__A2 _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_145_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_hold18_I net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10066_ _04661_ _04656_ _04662_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_4_4__f_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09720__A1 _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10011__I _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08287__B2 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _05401_ _05398_ _05402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10899_ as2650.chirpchar\[3\] _05256_ _05338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09787__A1 net210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__B _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_113_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_1595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06090_ net232 net251 _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_74_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_1568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07476__B _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08800_ as2650.stack\[15\]\[9\] _03495_ _02541_ as2650.stack\[14\]\[9\] _02520_ _03496_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_158_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09780_ _01526_ _04461_ _04462_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06992_ _01902_ _01756_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08731_ _01963_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05943_ _00740_ _00622_ _00589_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_1_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_68_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08514__A2 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09711__A1 _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09711__B2 _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08662_ _01789_ _01788_ _03270_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05874_ _00876_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_152_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07613_ _02390_ _02400_ _02402_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08593_ _01966_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_89_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07544_ wb_counter\[6\] _02346_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_92_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10856__I _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07475_ _02090_ wb_counter\[30\] _02273_ _02295_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09214_ _03895_ _03899_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_134_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06426_ net208 net191 net200 _01031_ _01185_ _01187_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__08326__I _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09227__B1 _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07230__I _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_62_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09145_ _03670_ _03671_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06357_ _01170_ _01171_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09778__B2 _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07789__B1 _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07789__C2 _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06288_ _00645_ _01128_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A1 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09076_ _03718_ _03764_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08027_ as2650.indirect_target\[5\] _02654_ _02780_ _02782_ _02783_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_13_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_57_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09950__A1 _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_89_wb_clk_i clknet_4_10__leaf_wb_clk_i clknet_leaf_89_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_21_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09978_ as2650.stack\[4\]\[3\] _04598_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_18_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_71_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08929_ _01211_ _01631_ _03620_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_77_1731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09106__B _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07405__I _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10822_ _01492_ net219 _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10753_ _05163_ _05215_ _05217_ _05218_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_54_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_153_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10684_ _05177_ _05175_ _05176_ _00795_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_168_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09769__A1 _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10379__A2 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05893__I3 _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11305_ _00101_ clknet_leaf_140_wb_clk_i net271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11236_ _00032_ clknet_leaf_117_wb_clk_i as2650.stack\[12\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09941__A1 _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11167_ _05467_ _05535_ _05540_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_8_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06755__A1 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10118_ _01083_ _04696_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_78_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11098_ _05436_ _05495_ _05498_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10049_ _04649_ _04646_ _04650_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06507__A1 _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05590_ as2650.indirect_target\[3\] _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_114_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_1762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05869__I0 _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07260_ _02090_ _02108_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07483__A2 net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08680__A1 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06211_ _01152_ _01169_ _01183_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_166_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07191_ _02035_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _01114_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold107_I wbs_dat_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06073_ _01053_ _01054_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_44_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09901_ as2650.cycle\[1\] _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_112_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09932__A1 _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09832_ _02568_ _04509_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_1842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06746__A1 _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10542__A2 _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ _02666_ _03065_ _04440_ _04443_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06975_ _01886_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08714_ as2650.stack\[12\]\[6\] _03411_ _03412_ as2650.stack\[13\]\[6\] _03413_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05926_ _00661_ _00804_ _00808_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_119_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09694_ as2650.cycle\[10\] _01528_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_59_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer10 _04059_ net354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07225__I _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09160__A2 _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ _03235_ _03322_ _03346_ _03234_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_96_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05857_ _00845_ as2650.regs\[1\]\[1\] _00864_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_90_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10845__A3 _05286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08576_ _03235_ _03236_ _03279_ _03234_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_33_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05788_ _00798_ net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_14_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07527_ wb_counter\[3\] _02327_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__09999__A1 _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_136_wb_clk_i clknet_4_3__leaf_wb_clk_i clknet_leaf_136_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_46_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07474__A2 _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ net284 _02282_ _02275_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08671__B2 _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06409_ _00857_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07389_ _02211_ wb_counter\[16\] _02223_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09128_ _01806_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output183_I net183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07226__A2 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_1465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06434__B1 _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _03706_ _03714_ _03719_ _03750_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__06985__A1 _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08187__B1 _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11021_ _01776_ _05445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_79_1826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_1363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08659__C _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05960__A2 _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_155_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07701__A3 _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_155_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11854_ net301 net180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_68_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08394__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ as2650.stack\[6\]\[12\] _05250_ _05251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11785_ _00564_ clknet_leaf_132_wb_clk_i as2650.stack\[13\]\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold85_I wbs_dat_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10736_ _05102_ _05202_ _05207_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10667_ _05164_ _05165_ _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_153_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_106_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10598_ as2650.stack\[7\]\[1\] _05118_ _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07738__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput108 net108 RAM_end_addr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput119 net119 RAM_end_addr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06976__A1 _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11219_ as2650.stack\[9\]\[15\] _05569_ _05573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10524__A2 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06760_ as2650.debug_psu\[2\] _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05711_ _00723_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06691_ _01044_ _01496_ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09693__A3 _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08430_ _03128_ _03149_ _02809_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05642_ _00654_ _00655_ _00591_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08361_ net207 _01437_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07312_ net135 _02139_ _02122_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_138_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_138_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08292_ _03018_ _03019_ _02622_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06259__A3 _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07243_ _02077_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_41_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07174_ net84 net116 _02041_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06125_ _01097_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_44_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06967__A1 _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06056_ _01038_ net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_61_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout302 net164 net302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09815_ _02473_ _03754_ _03573_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_96_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08184__A3 _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06195__A2 _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _02559_ _02568_ _02560_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_06958_ _01715_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05909_ _00914_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_96_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09677_ _04332_ _04355_ _04362_ _04354_ _03699_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_55_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_48_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _00694_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_48_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_312 io_oeb[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_70_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08628_ as2650.stack\[11\]\[3\] _03264_ _03290_ as2650.stack\[10\]\[3\] _03330_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xwrapped_as2650_323 la_data_out[44] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_334 la_data_out[37] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_167_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09170__I _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ as2650.stack\[12\]\[1\] _03261_ _03262_ as2650.stack\[13\]\[1\] _03263_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_132_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07447__A2 _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11570_ _00354_ clknet_leaf_127_wb_clk_i as2650.stack\[3\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10521_ _04653_ _05059_ _05064_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_1527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10452_ _04621_ _05019_ _05022_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10383_ _02781_ _04728_ _04761_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_wb_clk_i clknet_4_4__leaf_wb_clk_i clknet_leaf_33_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06034__I _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08389__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11004_ _05407_ _05430_ _05431_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_169_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_1412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08883__A1 _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05697__A1 _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11115__I _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07438__A2 _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11768_ _00547_ clknet_leaf_32_wb_clk_i as2650.stack\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08852__C _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10719_ as2650.stack\[8\]\[4\] _05197_ _05198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11699_ _00483_ clknet_leaf_14_wb_clk_i as2650.stack\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xrebuffer1 _00733_ net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_125_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09964__B _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09060__A1 _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10745__A2 _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07930_ _02677_ _02678_ _02656_ _02688_ _02689_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_122_1569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07861_ _01178_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_127_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09600_ _03728_ _04252_ _04278_ _04281_ _04285_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_0_39_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06812_ net188 _01732_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07792_ _02560_ _01513_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_88_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09531_ _03622_ _03639_ _03644_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_30_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06743_ _00662_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_30_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07931__C _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _04140_ _04115_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06674_ net254 _01602_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08413_ as2650.stack\[7\]\[15\] _02539_ _02542_ as2650.stack\[6\]\[15\] _03133_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05625_ as2650.indirect_target\[14\] _00635_ _00628_ as2650.page_reg\[1\] _00639_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_91_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09393_ _04076_ _04077_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_43_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08344_ _02553_ _03061_ _03062_ _03065_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_58_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08275_ _02997_ _03004_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07226_ wb_feedback_delay net105 _02005_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_104_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09051__A1 _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07157_ net76 net126 _02030_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06108_ as2650.warmup\[0\] as2650.warmup\[1\] net256 _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_4
X_07088_ _01869_ _01980_ _01985_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_37_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06039_ _01024_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_100_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05693__I _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output146_I net146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10104__I _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09729_ _03729_ _02585_ _03782_ _04413_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
Xclkbuf_leaf_151_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_151_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_69_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08865__A1 _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07413__I _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11622_ _00406_ clknet_leaf_24_wb_clk_i as2650.stack\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10774__I _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11553_ _00337_ clknet_leaf_41_wb_clk_i as2650.stack\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08093__A2 _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10504_ as2650.stack\[1\]\[4\] _05054_ _05055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08244__I _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11484_ _00268_ clknet_leaf_50_wb_clk_i as2650.irqs_latch\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10435_ _04393_ _04764_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_hold48_I net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09593__A2 _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10366_ _01387_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05603__A1 as2650.indirect_target\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05603__B2 as2650.PC\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06699__I _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10297_ _04842_ _04843_ _04873_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_97_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08553__B1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10014__I _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08847__C _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_83_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08856__A1 _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07323__I _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_1659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10663__A1 _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10663__B2 _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06390_ _01021_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_55_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06619__B1 _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10415__A1 _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08060_ _02813_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_12_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07011_ _01725_ _01920_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_1767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_77_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08792__B1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08962_ _03597_ _03652_ _03653_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_110_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ _01086_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_32_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08893_ _03584_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07198__I1 net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07844_ _01002_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_93_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07775_ _02524_ _02531_ _02538_ _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_75_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09514_ _04198_ _04199_ _03683_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_71_1704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06726_ _01640_ net347 _01650_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_91_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09445_ _04129_ _04130_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06657_ _01515_ _01583_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_91_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05608_ as2650.indirect_target\[8\] _00621_ _00615_ as2650.PC\[8\] _00622_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_168_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09376_ _03982_ _03987_ _03988_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06588_ _01526_ _01536_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__10406__A1 _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08327_ _03034_ _01299_ _03049_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_23_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10406__B2 _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10957__A2 _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ as2650.instruction_args_latch\[6\] _02975_ _02989_ _02981_ _02990_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07822__A2 _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07209_ net67 _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08189_ _02747_ _02931_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_132_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10709__A2 _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _04701_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_113_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10151_ _01237_ _01099_ _03727_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput280 net280 wbs_dat_o[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput291 net291 wbs_dat_o[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06312__I _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10082_ as2650.stack\[3\]\[3\] _04670_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_1499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_135_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07189__I1 net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_162_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07889__A2 _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08838__A1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10984_ _05404_ _05416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06313__A2 _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07510__A1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11605_ _00389_ clknet_leaf_6_wb_clk_i as2650.stack\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08066__A2 _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11536_ _00320_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11467_ _00251_ clknet_leaf_59_wb_clk_i as2650.debug_psl\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_169_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10418_ as2650.regs\[5\]\[7\] _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09566__A2 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11398_ _00182_ clknet_leaf_47_wb_clk_i as2650.indirect_target\[2\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08774__B1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10349_ _04918_ _04920_ _04923_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07329__A1 _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05890_ _00895_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10333__B1 _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10679__I _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06552__A2 _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07560_ wb_counter\[9\] _02359_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_152_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07053__I _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_100_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06511_ _01471_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_66_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09689__B _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07491_ web_behavior\[1\] _02305_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09230_ _03913_ _03915_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06442_ _01371_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06892__I _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09161_ _03823_ _03824_ _03847_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_100_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06373_ _01205_ _01207_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_20_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08112_ as2650.indirect_target\[10\] _01255_ _02848_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11061__A1 as2650.stack\[0\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09092_ _03780_ _03781_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08043_ _02796_ _02773_ _02797_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__09006__A1 _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ as2650.stack\[4\]\[9\] _04610_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07228__I _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08945_ _03623_ _03624_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05594__A3 _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08876_ as2650.stack\[8\]\[12\] _03516_ _03517_ as2650.stack\[9\]\[12\] _03464_ _03569_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05971__I _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input22_I bus_in_sid[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07827_ _01574_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08059__I _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07758_ _02526_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06709_ net248 net238 _01600_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07689_ net233 _01628_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output109_I net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08296__A2 _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__A1 _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09428_ _04100_ _04109_ _04113_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09359_ _01030_ _01021_ _04044_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_35_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09796__A2 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11321_ _00117_ clknet_leaf_139_wb_clk_i net289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_105_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11252_ _00048_ clknet_leaf_118_wb_clk_i as2650.stack\[11\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10273__B _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ _04781_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_164_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11183_ as2650.stack\[9\]\[0\] _05551_ _05552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10134_ _04711_ _04712_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06042__I _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10065_ as2650.stack\[10\]\[14\] _04657_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08397__C _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09720__A2 _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_158_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08287__A2 _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10967_ _04768_ _05399_ _05400_ _05401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06298__A1 _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_14_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10898_ net190 _04933_ _05304_ _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09236__A1 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06217__I _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08633__S _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_152_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11519_ _00303_ clknet_leaf_75_wb_clk_i as2650.ext_io_addr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_74_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06470__A1 _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06991_ _01901_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07970__A1 _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08730_ _01687_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_147_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05942_ _00944_ as2650.instruction_args_latch\[9\] _00945_ _00946_ _00947_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__06887__I _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09711__A2 _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08661_ _03356_ _03361_ _02550_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XANTENNA__08514__A3 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05873_ _00859_ _00876_ _00879_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_1_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07612_ net82 _02394_ _02401_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08592_ as2650.stack\[0\]\[2\] _03292_ _03293_ as2650.stack\[1\]\[2\] _03294_ _03295_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_152_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10609__A1 _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07543_ _02131_ wb_counter\[5\] _02336_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_76_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08278__A2 as2650.instruction_args_latch\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07474_ net111 _02119_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09213_ _03896_ _03897_ _03898_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_88_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06425_ _00910_ net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09227__A1 _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09227__B2 _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_1664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09144_ _03829_ _03830_ _03622_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__11034__A1 _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06356_ as2650.cycle\[11\] _01245_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06127__I _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07789__A1 net216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07789__B2 _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09075_ _01293_ _03764_ _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06287_ _01258_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_32_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08026_ _02781_ _02661_ _02741_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_4_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09950__A2 _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09977_ _01777_ _04596_ _04601_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08928_ _01768_ _01211_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output226_I net226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ _02871_ _03053_ _03552_ _03502_ _02736_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_77_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10821_ _05262_ _05263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_93_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ as2650.regs\[6\]\[0\] _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09122__B _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07421__I _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10683_ _04961_ _05177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_1450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_166_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11304_ _00100_ clknet_leaf_140_wb_clk_i net270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11235_ _00031_ clknet_leaf_116_wb_clk_i as2650.stack\[12\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06204__A1 net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11166_ as2650.stack\[13\]\[11\] _05536_ _05540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_8_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06755__A2 _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _01292_ _01243_ _03715_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_60_1791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11097_ as2650.stack\[14\]\[0\] _05497_ _05498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09083__I _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10048_ as2650.stack\[10\]\[9\] _04647_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_106_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06500__I _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold90 wbs_adr_i[19] net436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_89_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10022__I _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_63_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06210_ _01182_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_27_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06691__A1 _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07190_ _02050_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06141_ _00700_ _01110_ _01112_ _01113_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__08432__A2 _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06072_ _01052_ _00880_ _00858_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09900_ _04428_ _04553_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_93_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09831_ as2650.debug_psu\[7\] _02992_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06746__A2 _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06974_ as2650.debug_psu\[1\] _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09762_ _04438_ _04442_ _04445_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05925_ _00925_ _00929_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_08713_ _02494_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09693_ _02814_ _04373_ _04378_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11028__I _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer11 net256 net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08644_ _03194_ _03323_ _03345_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05856_ _00723_ _00863_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08575_ _02762_ _03239_ _03276_ _03278_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_117_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05787_ _00708_ _00795_ _00797_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09448__A1 net194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07526_ _02320_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07457_ _02078_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_146_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06682__A1 _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06408_ _00881_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07388_ _02212_ _02221_ _02222_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_66_1411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09127_ _03153_ _03811_ _03814_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06339_ _01307_ _01287_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_60_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07226__A3 _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_105_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_105_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_59_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09620__A1 _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09168__I _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06434__A1 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09058_ _03714_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08009_ _02765_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_41_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_83_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11020_ _05443_ _05439_ _05444_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09923__A2 _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_146_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06737__A2 _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11853_ net303 net163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_155_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10804_ _05231_ _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08247__I _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11784_ _00563_ clknet_leaf_25_wb_clk_i as2650.stack\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08111__A1 _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10735_ as2650.stack\[8\]\[11\] _05203_ _05207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06990__I _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10666_ _01808_ _04699_ _05165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_24_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10597_ _05071_ _05116_ _05119_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09611__A1 _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput109 net109 RAM_end_addr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_107_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08178__A1 _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11218_ _05475_ _05568_ _05572_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07925__A1 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11149_ _05523_ _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06230__I _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05710_ _00690_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_144_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10288__A2 _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06690_ net255 _01007_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08350__A1 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05641_ _00638_ _00639_ _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10687__I _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06900__A2 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08360_ _03077_ _03080_ _03081_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08157__I _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08102__A1 _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07061__I _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07311_ _02113_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_3_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_3_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08291_ _03007_ _02861_ _01256_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10835__I1 _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08653__A2 _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07242_ _02082_ _02089_ _02092_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_99_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07173_ _02035_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09602__A1 _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _01096_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_41_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06405__I net189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06055_ _01035_ _01037_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_169_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08169__A1 _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09905__A2 net147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout303 net164 net303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_39_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09814_ _04445_ _04478_ _04494_ _03534_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_35_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09745_ _01261_ _01324_ _01705_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_06957_ _01803_ _01869_ _01870_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_20_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_129_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05908_ _00913_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09676_ _04356_ _04357_ _04359_ _04361_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06888_ _01752_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_69_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08341__A1 _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_313 io_oeb[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_48_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ _03325_ _03326_ _03327_ _03328_ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05839_ as2650.regs\[2\]\[0\] _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xwrapped_as2650_324 la_data_out[45] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_335 la_data_out[38] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_90_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08558_ _03250_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_1481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07509_ _02317_ net411 _02318_ _02236_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_65_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08489_ _03193_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_108_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10520_ as2650.stack\[1\]\[11\] _05060_ _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07852__B1 _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output293_I net293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10451_ as2650.stack\[2\]\[0\] _05021_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10382_ _04940_ _04791_ _04951_ _04955_ _04826_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_81_1728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11003_ _05384_ _05396_ _05416_ as2650.regs\[0\]\[6\] _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_wb_clk_i clknet_4_15__leaf_wb_clk_i clknet_leaf_73_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08332__A1 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08883__A2 _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06894__A1 _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11767_ _00546_ clknet_leaf_32_wb_clk_i as2650.stack\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_4_14__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10718_ _05190_ _05197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_99_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11698_ _00482_ clknet_leaf_99_wb_clk_i as2650.regs\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_133_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10649_ as2650.regs\[1\]\[2\] _05154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xrebuffer2 net345 net346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09899__A1 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09899__B2 as2650.trap vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ _02623_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07056__I _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06811_ _01730_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_120_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07791_ _01459_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_39_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06742_ net245 _01602_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09530_ _02469_ _04211_ _04213_ _04215_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_30_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06895__I as2650.PC\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09461_ _04135_ _04139_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06673_ _01006_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10130__A1 _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05624_ _00633_ _00637_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05688__A2 _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08412_ as2650.stack\[0\]\[15\] _02527_ _02530_ as2650.stack\[1\]\[15\] _03131_ _03132_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_4_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09392_ _04076_ _04077_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_0_87_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_43_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08343_ _03064_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08626__A2 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09823__A1 net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _02998_ _02637_ _02999_ _01259_ _03003_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_46_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07225_ _02076_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11041__I _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07156_ _02031_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09051__A2 _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10197__A1 _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06107_ _01080_ net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_112_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07087_ as2650.stack\[11\]\[7\] _01981_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input52_I ram_bus_in[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06038_ _01023_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_1768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_125_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08011__B1 _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_137_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08562__A1 _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output139_I net139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07989_ as2650.ivectors_base\[0\] _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_74_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _04186_ _04412_ _04193_ _03724_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09659_ _02715_ _01632_ _01643_ _02726_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10121__A1 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11621_ _00405_ clknet_leaf_18_wb_clk_i as2650.stack\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_120_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_120_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_166_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_146_Left_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06628__A1 _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11552_ _00336_ clknet_leaf_41_wb_clk_i as2650.stack\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10503_ _05047_ _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11483_ _00267_ clknet_leaf_51_wb_clk_i as2650.irqs_latch\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10434_ _01085_ _04426_ _05001_ _05005_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10188__A1 _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10365_ as2650.regs\[5\]\[5\] _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_123_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08260__I _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10296_ _04844_ _04872_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_155_Left_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_1581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07356__A2 _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_70_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10360__A1 _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07108__A2 _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08305__B2 net208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11126__I _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06867__A1 _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10030__I _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_164_Left_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09805__A1 _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06619__A1 wb_debug_cc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10966__A3 _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07010_ _01919_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09569__B1 _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07044__A1 net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08961_ _03594_ _03596_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_99_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07912_ _02668_ _02671_ _02672_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08892_ _03583_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_32_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07843_ _02449_ _02609_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_120_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10351__A1 _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06839__B _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07774_ as2650.stack\[15\]\[13\] _02539_ _02542_ as2650.stack\[14\]\[13\] _02521_
+ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07514__I _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09513_ _03607_ _03647_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06725_ _01640_ _01031_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08847__A2 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09444_ _04108_ _04124_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06656_ _01589_ _01590_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_166_Right_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05607_ _00599_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06587_ net237 _01527_ _01531_ _01535_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_136_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09375_ _04060_ _04053_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_148_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08326_ _01330_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08345__I _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08257_ _02968_ _02987_ _02988_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07208_ _01119_ _02059_ _02061_ _02063_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_105_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08188_ _01293_ _01306_ _02930_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_104_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07139_ net99 net133 _02020_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08783__A1 _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10150_ _04705_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_1445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output256_I net355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput270 net270 wbs_dat_o[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput281 net281 wbs_dat_o[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_101_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput292 net292 wbs_dat_o[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10081_ _04631_ _04668_ _04673_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09904__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10342__A1 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06010__A2 _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10983_ _05317_ _05409_ _05414_ _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_38_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11604_ _00388_ clknet_leaf_10_wb_clk_i as2650.stack\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06077__A2 net248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11535_ _00319_ clknet_leaf_16_wb_clk_i as2650.stack\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold60_I net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09015__A2 _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11466_ _00250_ clknet_leaf_60_wb_clk_i as2650.debug_psl\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08223__B1 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10417_ _04967_ _04787_ _04986_ _04724_ _04989_ _04771_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_11397_ _00181_ clknet_leaf_49_wb_clk_i as2650.indirect_target\[1\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09086__I _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06503__I _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10348_ _04921_ _04922_ _04882_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_72_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10025__I _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10279_ _04853_ _04855_ _04742_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07329__A2 _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08526__B2 _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07762__C _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07334__I _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_1451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08829__A2 _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05760__A1 _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06510_ _01260_ _01267_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07490_ _02057_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_66_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06441_ _01390_ _01339_ _01398_ _01399_ _01403_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_29_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_5_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05789__I net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09160_ _03607_ _03776_ _03837_ _03846_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_25_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06372_ _01287_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_25_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_100_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09254__A2 _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08111_ _02861_ _02740_ _02741_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_44_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09091_ _03657_ _03776_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11061__A2 _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08042_ _01160_ _01829_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07937__C _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07017__A1 _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05579__A1 as2650.relative_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09993_ _01883_ _04609_ _04611_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _03632_ _03634_ _03635_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08768__C _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08875_ as2650.stack\[11\]\[12\] _03495_ _02541_ as2650.stack\[10\]\[12\] _03568_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07826_ _02463_ _02594_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07244__I _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I bus_in_serial_ports[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07757_ _02525_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_75_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06708_ _01628_ _01634_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10627__A2 _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07688_ net252 net238 _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ _04110_ _04111_ _04112_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_149_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06639_ _01575_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09358_ _04010_ _04011_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08309_ _03034_ as2650.instruction_args_latch\[12\] _03026_ _03035_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07256__A1 _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09289_ _03959_ _03960_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11320_ _00116_ clknet_leaf_102_wb_clk_i net287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_69_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11251_ _00047_ clknet_leaf_119_wb_clk_i as2650.stack\[11\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10202_ _01697_ _04183_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_24_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11182_ _05550_ _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_164_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _01461_ _01483_ _04701_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_98_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10064_ _01953_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10315__A1 _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__A1 _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07154__I _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1057 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10966_ _03817_ as2650.regs\[4\]\[0\] _01547_ _05400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_116_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10897_ _03335_ _05321_ _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_14_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_117_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09236__A2 _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11518_ _00302_ clknet_leaf_54_wb_clk_i net145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08713__I _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06470__A2 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11449_ _00233_ clknet_leaf_32_wb_clk_i as2650.ivectors_base\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08747__A1 _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06990_ _01682_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input7_I bus_in_gpios[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ _00589_ _00940_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09172__A1 _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09172__B2 _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_1693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05872_ _00657_ _00877_ _00878_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_1_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08660_ _03357_ _03358_ _03359_ _03360_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_1_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07611_ _02384_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_163_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05733__A1 _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08591_ _02503_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_152_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07542_ _02341_ _02343_ _02345_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_152_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__A1 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07473_ _02277_ _02291_ _02294_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08683__B1 _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11461__D _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09212_ _00717_ _01498_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06424_ _01347_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06408__I _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07238__A1 _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09143_ _03625_ _03666_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06355_ _01319_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09074_ _02919_ _02586_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_44_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06286_ _01257_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_142_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08025_ _02770_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_130_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07239__I _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_57_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10545__A1 _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09976_ as2650.stack\[4\]\[2\] _04598_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08927_ _03617_ _03618_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05972__A1 _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08858_ _03190_ _01920_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_38_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08910__A1 _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output121_I net121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07809_ _01188_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output219_I net219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08789_ _01879_ _03459_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10820_ _05255_ _05262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_wb_clk_i clknet_4_11__leaf_wb_clk_i clknet_leaf_98_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10751_ _05216_ _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_82_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _05174_ _05175_ _05176_ _00916_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_153_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07858__B _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11025__A2 _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_166_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11303_ _00099_ clknet_leaf_141_wb_clk_i net269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08729__A1 _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11234_ _00030_ clknet_leaf_117_wb_clk_i as2650.stack\[12\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_1771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11165_ _05465_ _05535_ _05539_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10116_ _04693_ _04694_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11096_ _05496_ _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08201__C _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09154__A1 _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10047_ _01898_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10839__A2 _05279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold80 net458 net424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__08901__A1 _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold91 _02068_ net437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_0_118_1553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09701__I0 net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07468__A1 net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10949_ as2650.regs\[4\]\[6\] _05335_ _05384_ _05294_ _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08665__B1 _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__I2 net196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08871__C _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11016__A2 _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06691__A2 _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06140_ as2650.insin\[2\] _00700_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08968__A1 _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08443__I _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10775__A1 as2650.stack\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_1660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08432__A3 _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06071_ _01052_ _00858_ _00880_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_129_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07059__I _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08196__A2 _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09830_ net37 _02480_ _04507_ _02483_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_123_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09761_ _04444_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05954__A1 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06973_ _01871_ _01883_ _01885_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11456__D _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08712_ _02487_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05924_ _00811_ _00927_ _00928_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10213__I _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09692_ _02766_ _02791_ _02781_ _04377_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_94_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xrebuffer12 _01357_ net356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08643_ _03225_ _03340_ _03342_ _03344_ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_55_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05855_ as2650.regs\[5\]\[1\] _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08574_ _03277_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05786_ _00796_ as2650.regs\[6\]\[5\] _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09448__A2 _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07525_ _02321_ _02329_ _02331_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08656__B1 _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06138__I _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07456_ _02278_ wb_counter\[26\] _02273_ _02280_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_46_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06407_ _01368_ _01369_ _01370_ _00895_ _01185_ _01187_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_161_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07387_ _02183_ _01565_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_1495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09126_ _03813_ _03757_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06338_ _01098_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_59_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06269_ _01240_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_115_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09057_ net188 _03723_ _03740_ _03748_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08008_ net62 _02763_ _02764_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_104_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_145_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_145_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_143_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__A2 _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06601__I _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09959_ net224 _04586_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11852_ net302 net162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_155_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_155_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10803_ _05229_ _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_67_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11783_ _00562_ clknet_leaf_24_wb_clk_i as2650.stack\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08972__B _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_4_13__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10734_ _05100_ _05202_ _05206_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10793__I _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10665_ _04714_ _04720_ _04307_ _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_84_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10596_ as2650.stack\[7\]\[0\] _05118_ _05119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09611__A2 _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_131_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11217_ as2650.stack\[9\]\[14\] _05569_ _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07925__A2 _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11148_ _05521_ _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_78_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09127__A1 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10033__I _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11079_ _05172_ _05480_ _05482_ _05485_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__09822__I _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05640_ _00652_ _00647_ _00653_ _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _02130_ _02153_ _02154_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08290_ _02997_ _03017_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07161__I0 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07241_ _02090_ _02091_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_99_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_99_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07172_ _02040_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_hold112_I wbs_dat_i[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06123_ _01095_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06054_ _00770_ _01036_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_125_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08169__A2 _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_115_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09813_ _02748_ _04482_ _04493_ _04444_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_35_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09744_ _01087_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06956_ as2650.stack\[12\]\[7\] _01821_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08776__C _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05907_ _00912_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_74_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09675_ _04360_ _02731_ _02770_ _04282_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08877__B1 _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06887_ _00923_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_97_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08341__A2 _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_1758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08626_ as2650.stack\[4\]\[3\] _03305_ _03306_ as2650.stack\[5\]\[3\] _03298_ _03328_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_48_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_314 io_oeb[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_05838_ _00723_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_136_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06352__A1 _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_325 la_data_out[46] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_336 la_data_out[39] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_90_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08557_ _03248_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08629__B1 _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05769_ _00779_ _00617_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ net96 net437 _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08488_ _03190_ _03192_ _02655_ _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_108_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07152__I0 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10987__A1 _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07439_ _02064_ net120 _02011_ as2650.debug_psu\[7\] _02146_ _02266_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__07852__B2 _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_154_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ _05020_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output286_I net286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09109_ _01292_ _01294_ _01513_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_21_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10381_ _04756_ _04954_ _04882_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_115_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05615__B1 _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07907__A2 _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11002_ _05375_ _05403_ _05429_ _05430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09109__A1 _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08332__A2 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_42_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_42_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_169_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11219__A2 _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_hold90_I wbs_adr_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11766_ _00545_ clknet_leaf_26_wb_clk_i as2650.stack\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_81_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07143__I0 net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07843__A1 _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10717_ _05188_ _05196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_71_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11697_ _00481_ clknet_leaf_99_wb_clk_i as2650.regs\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_133_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10648_ _04834_ _05146_ _05149_ _04839_ _05151_ _05153_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
Xrebuffer3 _00924_ net347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10028__I _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10579_ _05075_ _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_90_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11155__A1 _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09899__A2 _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08020__A1 _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__I _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06810_ _01730_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08571__A2 _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07790_ _02466_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_159_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_88_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08596__C _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06741_ _01418_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08323__A2 _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09520__A1 _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09460_ _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06672_ _01600_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_133_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08168__I as2650.instruction_args_latch\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06334__A1 _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08411_ _03130_ _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05623_ _00634_ _00597_ _00636_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_1499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05688__A3 _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06885__A2 _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09391_ _04002_ _04003_ _03991_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_0_87_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08342_ _03063_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_43_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07134__I0 net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09823__A2 _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08273_ _03000_ _02603_ net204 _03002_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_50_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07224_ _02075_ wb_feedback_delay _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_67_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09587__A1 _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07155_ net75 net125 _02030_ _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09051__A3 _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06106_ _01079_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07086_ _01853_ _01980_ _01984_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_1459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06037_ _01022_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_1762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input45_I irqs[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07988_ _02720_ _02722_ _02743_ _02744_ _02745_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_57_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09727_ _04183_ _04156_ _04410_ _04411_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06939_ as2650.stack\[12\]\[6\] _01821_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09658_ _02715_ _01632_ _01621_ _02675_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_85_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output201_I net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08609_ _03058_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09589_ _04263_ _04259_ _04273_ _04274_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_11620_ _00404_ clknet_leaf_17_wb_clk_i as2650.stack\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08078__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06628__A2 _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11551_ _00335_ clknet_leaf_12_wb_clk_i as2650.stack\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _05045_ _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11482_ _00266_ clknet_leaf_50_wb_clk_i as2650.irqs_latch\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08742__S _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10433_ _04727_ _05004_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08541__I _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10364_ _04909_ _04789_ _04931_ _04835_ _04938_ _04840_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XANTENNA__08250__B2 net201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10295_ _04385_ _04846_ _04870_ _04871_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_104_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06061__I _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08697__B _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08553__A2 _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09750__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08305__A2 _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09502__A1 _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10112__A2 _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06867__A2 _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08069__A1 as2650.indirect_target\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07816__A1 _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06619__A2 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11749_ _00002_ clknet_leaf_88_wb_clk_i as2650.chirpchar\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09569__A1 _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_12_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08451__I _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08792__A2 _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08960_ _03604_ _03649_ _03651_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_45_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ as2650.wb_hidden_rom_enable _01538_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08891_ _01114_ _01209_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XTAP_TAPCELL_ROW_32_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07842_ as2650.insin\[1\] _02596_ _02600_ _02608_ _02604_ _02609_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_75_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07773_ _02541_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11464__D _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09512_ _03834_ _03835_ _03824_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06724_ net243 _01602_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09443_ _04121_ _04122_ _04120_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06655_ _01584_ _00179_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05606_ _00601_ _00619_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09374_ _03993_ _03996_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06586_ _01000_ _01255_ _01533_ _01534_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08325_ _03029_ _03047_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_1740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11052__I _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08256_ as2650.instruction_args_latch\[6\] _02978_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08480__A1 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ _02062_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08187_ _01998_ _01722_ _02653_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_127_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07138_ _02021_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07069_ _01971_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xoutput260 net260 rom_bus_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__11119__A1 as2650.stack\[14\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput271 net271 wbs_dat_o[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10590__A2 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output151_I net151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput282 net282 wbs_dat_o[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_100_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput293 net293 wbs_dat_o[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10080_ as2650.stack\[3\]\[2\] _04670_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_1588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output249_I net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09732__A1 _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10342__A2 _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07705__I _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10982_ _03813_ as2650.regs\[4\]\[2\] _03104_ _05414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_151_1531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11603_ _00387_ clknet_leaf_7_wb_clk_i as2650.stack\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11534_ _00318_ clknet_leaf_15_wb_clk_i as2650.stack\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11070__A3 _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_115_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11465_ _00249_ clknet_4_12__leaf_wb_clk_i as2650.debug_psl\[0\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08223__A1 _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _04157_ _04779_ _04988_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_111_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11396_ _00180_ clknet_leaf_122_wb_clk_i as2650.chirp_ptr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_111_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08774__A2 _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10347_ _03858_ _04819_ _04814_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10306__I _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10581__A2 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10278_ _01625_ _04854_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_104_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06388__I1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_1739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11137__I _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05760__A2 _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06440_ _01400_ _01402_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_111_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08446__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06371_ _01117_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_57_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08110_ as2650.instruction_args_latch\[10\] _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09090_ _01200_ _03695_ _03770_ _03779_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_160_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08041_ _02769_ _01829_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07017__A2 _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09962__A1 _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ as2650.stack\[4\]\[8\] _04610_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08943_ _03631_ _03628_ _03630_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_23_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08874_ _03563_ _03564_ _03565_ _03566_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06528__A1 _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07825_ _02481_ _02571_ _02593_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ _02489_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06707_ _01629_ _01633_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07687_ _01067_ _01552_ _02451_ _02458_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_39_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08150__B1 _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09426_ _00730_ _00793_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06638_ _01277_ _01152_ _01282_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_113_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09357_ _04032_ _04041_ _04042_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06569_ _01517_ _01519_ _01521_ net155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_164_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _03006_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_118_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07256__A2 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08453__A1 _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ _03965_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_output199_I net199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10260__A1 _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08239_ _02949_ _02973_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11250_ _00046_ clknet_leaf_121_wb_clk_i as2650.stack\[11\]\[13\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08205__A1 net213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10201_ _03658_ _04774_ _04776_ _04779_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_113_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11181_ _05547_ _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_164_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09915__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10132_ _01461_ _04701_ _04710_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_98_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09705__A1 _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10063_ _04659_ _04656_ _04660_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_1395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05990__A2 net255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__A2 _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_104_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10965_ _05143_ _05283_ _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_104_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_1609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10896_ _05287_ _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_156_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_113_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11517_ _00301_ clknet_leaf_54_wb_clk_i net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_113_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11448_ _00232_ clknet_leaf_33_wb_clk_i as2650.ivectors_base\[8\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09944__A1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08747__A2 _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10036__I _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11379_ _00175_ clknet_leaf_62_wb_clk_i as2650.insin\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06758__A1 net253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05940_ _00740_ _00622_ _00624_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_59_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05871_ _00588_ as2650.instruction_args_latch\[1\] _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_1_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07610_ wb_counter\[19\] _02399_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_50_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08590_ _02497_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_117_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05733__A2 as2650.instruction_args_latch\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07541_ net362 _02344_ _02330_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07472_ net287 _02282_ _02293_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07080__I _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09211_ _00755_ _00824_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06423_ _00805_ _01340_ _01341_ _01384_ _01386_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09142_ _03827_ _03828_ _03627_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_72_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06354_ _01318_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08435__A1 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__A2 _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10242__A1 _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08986__A2 _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09073_ _03752_ _03763_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06285_ _01253_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08024_ _02698_ _02779_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06749__A1 _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10545__A2 _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__C _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09975_ _01760_ _04596_ _04600_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08926_ _02613_ _03584_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_1569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08857_ _02935_ _01915_ _03550_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07808_ _02576_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08910__A2 _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08788_ _01893_ _03351_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05724__A2 _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07739_ _01689_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output114_I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10750_ _05168_ _05214_ _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_157_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_4_12__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09409_ _00758_ _01030_ _00827_ _00720_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_95_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10681_ _05169_ _05176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_165_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_wb_clk_i clknet_4_13__leaf_wb_clk_i clknet_leaf_67_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11302_ _00098_ clknet_leaf_143_wb_clk_i net268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08729__A2 _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11233_ _00029_ clknet_leaf_126_wb_clk_i as2650.stack\[12\]\[12\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11164_ as2650.stack\[13\]\[10\] _05536_ _05539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10115_ _01727_ _01697_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11095_ _05493_ _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_159_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09154__A2 _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10046_ _04645_ _04646_ _04648_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_106_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold70 net453 net414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_76_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold81 net467 net425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold92 wbs_dat_i[29] net438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09701__I1 net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10948_ _04322_ _05280_ _05383_ _05384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08665__A1 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08665__B2 _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05869__I3 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10879_ as2650.regs\[4\]\[2\] _05288_ _05319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10224__B2 _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09090__A1 _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__A1 as2650.PC\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06070_ _01043_ _00881_ _00879_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_1 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07640__A2 wb_counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05651__A1 as2650.wb_hidden_rom_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_105_wb_clk_i_I clknet_4_8__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10527__A2 _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09760_ _04443_ _02666_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06972_ as2650.stack\[12\]\[8\] _01884_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ as2650.stack\[8\]\[6\] _02488_ _02495_ as2650.stack\[9\]\[6\] _02501_ _03410_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05923_ _00811_ as2650.instruction_args_latch\[4\] _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09691_ _02607_ _02640_ _02616_ _02619_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_98_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08642_ _03343_ _02655_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xrebuffer13 _00938_ net429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
X_05854_ _00847_ _00860_ _00861_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08573_ _03230_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_132_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05785_ _00724_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07524_ net94 _02323_ _02330_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08656__B2 as2650.stack\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07455_ net107 _02279_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_9_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_46_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06406_ net197 _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07386_ net106 _02199_ _02213_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_144_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09125_ _03812_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06337_ _01305_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_45_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11060__I _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09056_ _03733_ _03746_ _03747_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06268_ _01239_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_108_1745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08007_ _02763_ _01176_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_1756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06199_ _01170_ _01171_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_130_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__B1 _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09958_ _01488_ _01639_ _04589_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_102_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05945__A2 as2650.instruction_args_latch\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output231_I net231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08909_ _03586_ _01660_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_142_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_114_wb_clk_i clknet_4_10__leaf_wb_clk_i clknet_leaf_114_wb_clk_i vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09889_ as2650.stack\[5\]\[12\] _04546_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_159_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11851_ net302 net170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_155_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_1749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10802_ _05102_ _05243_ _05248_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06329__I _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08647__A1 _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11782_ _00561_ clknet_leaf_26_wb_clk_i as2650.stack\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10733_ as2650.stack\[8\]\[10\] _05203_ _05206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08544__I _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10664_ _04768_ _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ _05117_ _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_69_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09072__B2 _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09611__A3 _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_1844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11216_ _05473_ _05568_ _05571_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08178__A3 _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06189__A2 _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07386__A1 net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11147_ _05447_ _05522_ _05528_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05936__A2 _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11078_ as2650.regs\[7\]\[2\] _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_159_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10029_ _04624_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_76_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07161__I1 net128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07240_ wb_counter\[0\] _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_99_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07171_ net82 net115 _02036_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06122_ _00700_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold105_I wbs_dat_i[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06053_ _00784_ _00810_ net348 _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_61_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09812_ _02599_ _04489_ _04492_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_1653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06955_ _01868_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09743_ _04424_ _04426_ _04427_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05906_ as2650.regs\[1\]\[4\] as2650.regs\[5\]\[4\] _00789_ _00912_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_154_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09674_ _01401_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06886_ _01715_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08625_ as2650.stack\[7\]\[3\] _03264_ _03290_ as2650.stack\[6\]\[3\] _03327_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_48_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05837_ as2650.regs\[1\]\[0\] as2650.regs\[5\]\[0\] _00845_ _00846_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_315 io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_90_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11055__I _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_326 la_data_out[47] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_6_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xwrapped_as2650_337 la_data_out[40] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_08556_ as2650.stack\[8\]\[1\] _03249_ _03251_ as2650.stack\[9\]\[1\] _03252_ _03260_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05768_ _00613_ _00616_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07507_ as2650.wb_hidden_rom_enable _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08792__C _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _03191_ _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05699_ _00712_ net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_65_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07152__I1 net124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07438_ _02251_ _02264_ _02265_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09054__A1 _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ net127 _02199_ _02175_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09054__B2 _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10739__A2 _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09108_ _03767_ _03793_ _03797_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _01657_ _04818_ _04953_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_output181_I net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_148_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05615__B2 as2650.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09039_ _03730_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_60_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11001_ _05428_ _01534_ _05403_ _05429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__07907__A3 _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08868__A1 _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08332__A3 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06059__I _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10427__A1 _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11765_ _00544_ clknet_leaf_25_wb_clk_i as2650.stack\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_81_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_82_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_82_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07143__I1 net135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_hold83_I _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10716_ _05082_ _05189_ _05195_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11696_ _00480_ clknet_leaf_97_wb_clk_i as2650.regs\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_11_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05854__A1 _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10647_ as2650.regs\[1\]\[1\] _05153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_133_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer4 _00934_ net348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_94_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10578_ _05073_ _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05606__A1 _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08556__B1 _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10044__I _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10979__I _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06740_ _01657_ _01601_ _01663_ net171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_88_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08859__B2 _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10666__A1 _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06671_ _01531_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08410_ _02503_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_87_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05622_ as2650.indirect_target\[13\] _00635_ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _04073_ _04074_ _04075_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08341_ _01452_ _01475_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08087__A2 _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07134__I1 net131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08272_ _03001_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_62_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07223_ _02074_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05845__A1 _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07154_ _02014_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09587__A2 _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06105_ _00666_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07085_ as2650.stack\[11\]\[6\] _01981_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06036_ _00803_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_100_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08011__A2 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input38_I io_in[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07987_ _02673_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_138_1535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06938_ _01852_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09726_ _02477_ _03440_ _04189_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10657__A1 _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09657_ _02645_ _01608_ _01632_ _02715_ _01621_ _02675_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_39_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10657__B2 _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06869_ _01786_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_97_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08608_ _03300_ _03310_ _02550_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_96_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09588_ _01837_ _03856_ _04253_ _04254_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08539_ _01443_ _03057_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08078__A2 _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11550_ _00334_ clknet_leaf_12_wb_clk_i as2650.stack\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10501_ _04633_ _05046_ _05052_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11481_ _00265_ clknet_leaf_51_wb_clk_i as2650.irqs_latch\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09027__A1 _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10432_ _01674_ _04864_ _05003_ _04750_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_145_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _04936_ _04937_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_81_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08250__A2 _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06261__A1 _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10294_ _02716_ _04826_ _04845_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_70_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_69_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08269__I as2650.instruction_args_latch\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__I _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10648__A1 _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09502__A2 _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10648__B2 _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_83_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07816__A2 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11748_ _00001_ clknet_leaf_88_wb_clk_i as2650.chirpchar\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_78_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10039__I _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__A1 _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11679_ _00463_ clknet_leaf_23_wb_clk_i as2650.stack\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09569__A2 _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06252__I _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_36_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07910_ as2650.cpu_hidden_rom_enable _02670_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08890_ _02812_ _01213_ _03581_ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_166_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_32_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10887__A1 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _02607_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_87_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06555__A2 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10502__I _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _02540_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_100_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06723_ _01388_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09511_ _04184_ _04186_ _04192_ _04193_ _04196_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__07504__A1 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09442_ _03928_ _04089_ _04125_ _04127_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06654_ _00178_ _00179_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_133_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07811__I _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05605_ _00613_ _00616_ _00617_ _00618_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09373_ _04012_ _04016_ _04058_ _04046_ _04055_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__09257__A1 _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06585_ _01085_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08324_ _02761_ _03045_ _03046_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__C _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_30_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08255_ _02969_ _02803_ _02976_ net202 _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_117_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09009__A1 _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08480__A2 _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07206_ net66 _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08186_ _01269_ _01320_ _01334_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08768__B1 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ net98 net132 _02020_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07068_ _01972_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput250 net250 requested_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput261 net261 rom_bus_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput272 net272 wbs_dat_o[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06019_ _00914_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_11_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput283 net283 wbs_dat_o[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput294 net294 wbs_dat_o[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07194__S _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output144_I net144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10342__A3 _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09709_ _02670_ _04381_ _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_10981_ _05408_ _05411_ _05413_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_139_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07721__I _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11602_ _00386_ clknet_leaf_10_wb_clk_i as2650.stack\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06337__I _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire300 net185 net300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_65_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10802__A1 _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10263__C1 _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11533_ _00317_ clknet_leaf_2_wb_clk_i as2650.stack\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11464_ _00248_ clknet_leaf_43_wb_clk_i as2650.PC\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10415_ _01838_ _04932_ _04987_ _04964_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_104_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08223__A2 _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11395_ _00179_ clknet_leaf_29_wb_clk_i as2650.chirp_ptr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_111_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10346_ _02894_ _01393_ _04865_ _01395_ _04864_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_123_1623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold46_I net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_128_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06785__A2 _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10277_ as2650.debug_psl\[5\] _01614_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_124_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_1486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06370_ _01334_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_25_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08040_ _02786_ _01845_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_72_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09991_ _04597_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_1607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05579__A3 as2650.cycle\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08942_ _03633_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_99_1629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08873_ as2650.stack\[4\]\[12\] _02526_ _02529_ as2650.stack\[5\]\[12\] _03520_ _03566_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__11475__D _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07824_ _02573_ _02592_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ as2650.stack\[11\]\[13\] _01693_ _01969_ as2650.stack\[10\]\[13\] _02524_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06706_ _01604_ _01632_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07686_ net232 _02452_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_4_7__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09425_ _00720_ _01024_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06637_ _01573_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_133_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11063__I _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11037__A1 _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06157__I _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06568_ _01520_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09356_ _04017_ _04024_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_168_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_139_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_139_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08307_ _03029_ _03032_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09287_ _03963_ _03964_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09650__A1 _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06499_ _01151_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_117_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_1444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ as2650.instruction_args_latch\[3\] _02950_ _02972_ _02958_ _02973_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_117_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06464__A1 _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_1622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08169_ _02913_ _00652_ _01296_ _01722_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_82_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10200_ _04778_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_82_1655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06216__A1 _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11180_ _05548_ _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_164_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10131_ _01262_ _01297_ _01318_ _01471_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_105_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_164_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_1829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09705__A2 _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ as2650.stack\[10\]\[13\] _04657_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10964_ _05397_ _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_104_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10895_ _05333_ _05297_ _05298_ _00822_ _05334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_6_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__A2 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11516_ _00300_ clknet_leaf_53_wb_clk_i net143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11447_ _00231_ clknet_leaf_38_wb_clk_i as2650.ivectors_base\[7\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11200__A1 _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11378_ _00174_ clknet_leaf_62_wb_clk_i as2650.insin\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07955__A1 _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10329_ _03548_ _04775_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11148__I _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05870_ net305 _00836_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_94_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08885__C _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07540_ _02322_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_89_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07471_ _02292_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09880__A1 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__A2 _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06422_ _01367_ _01385_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09210_ _00791_ _01028_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ _03661_ _03628_ _03630_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_leaf_134_wb_clk_i_I clknet_4_2__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06353_ _01170_ _01317_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_169_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10242__A2 _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09072_ _03753_ _03759_ _03762_ _01295_ _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06284_ _01255_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_128_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08023_ as2650.indirect_target\[5\] _02635_ _02778_ _02708_ _02779_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_13_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08199__A1 _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07964__C _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_1415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09974_ as2650.stack\[4\]\[1\] _04598_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07536__I _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08925_ _01349_ _01225_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08856_ _01275_ _03537_ _03549_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input20_I bus_in_sid[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08371__A1 net212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07807_ _02575_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_05999_ as2650.cycle\[2\] as2650.cycle\[8\] _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08787_ _02636_ _03223_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07738_ as2650.stack\[0\]\[13\] _02493_ _02500_ as2650.stack\[1\]\[13\] _02506_ _02507_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08123__A1 as2650.instruction_args_latch\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output107_I net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07669_ wb_counter\[31\] _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_71_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_157_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06685__A1 _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09408_ _00730_ _01012_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10680_ _05166_ _05175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10481__A2 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09339_ _04017_ _04024_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09623__A1 _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11301_ _00097_ clknet_leaf_143_wb_clk_i net267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11232_ _00028_ clknet_leaf_135_wb_clk_i as2650.stack\[12\]\[11\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11163_ _05463_ _05535_ _05538_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_1458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_36_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_1795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10114_ _01228_ _03151_ _04432_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11094_ _05494_ _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_8_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10045_ as2650.stack\[10\]\[8\] _04647_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_106_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08362__A1 _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold60 net103 net404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold71 net439 net415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold82 wbs_cyc_i net426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold93 wbs_dat_i[27] net439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08114__A1 as2650.ivectors_base\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_1543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_63_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09701__I2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10947_ _05320_ _05382_ _05383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_128_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09862__A1 _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10878_ _05317_ _05284_ _05285_ _00894_ _05318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_155_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__A2 _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10047__I _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_2 _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09917__A2 _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07928__B2 _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06971_ _01738_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_52_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08710_ as2650.stack\[11\]\[6\] _01688_ _01964_ as2650.stack\[10\]\[6\] _03409_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05922_ _00779_ _00926_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09690_ _04373_ _04375_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_119_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08353__A1 net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05805__S _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08641_ _03190_ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_05853_ _00724_ as2650.regs\[7\]\[1\] _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xrebuffer14 _00619_ net430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_55_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08572_ _02685_ _03108_ _03240_ _03238_ _03275_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05784_ as2650.regs\[2\]\[5\] _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_1621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07523_ _02292_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_18_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08656__A2 _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07454_ _02245_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_1806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_46_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06405_ net189 _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_07385_ _02190_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_169_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09605__A1 _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06336_ _01304_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09124_ _01807_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09700__S1 _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09081__A2 _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07092__A1 _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09055_ _03721_ _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_5_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06267_ _01238_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_66_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08006_ _01153_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_143_1637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07219__I0 net161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09908__A2 _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06198_ _01127_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07919__A1 _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07266__I _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_146_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09957_ net223 _01545_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_5_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08908_ _03598_ _03599_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_77_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ _04527_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08344__A1 _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output224_I net224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08839_ _02673_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_169_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11850_ net302 net169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_101_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_154_wb_clk_i clknet_4_0__leaf_wb_clk_i clknet_leaf_154_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_16_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10801_ as2650.stack\[6\]\[11\] _05244_ _05248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_155_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08647__A2 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11781_ _00560_ clknet_leaf_25_wb_clk_i as2650.stack\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10732_ _05098_ _05202_ _05205_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10663_ _05011_ _05156_ _05157_ _05015_ _05158_ _05162_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_49_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10594_ _05114_ _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09611__A4 _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11215_ as2650.stack\[9\]\[13\] _05569_ _05571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_92_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08583__A1 _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06080__I net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11146_ as2650.stack\[13\]\[3\] _05524_ _05528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11077_ _05171_ _05480_ _05482_ _05484_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08335__A1 _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _01819_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_95_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06897__A1 _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09835__A1 _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__A2 _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_46_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10996__A3 _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_99_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_99_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07170_ _02039_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_41_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06121_ _01093_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07074__A1 _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10748__A3 _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06052_ _00982_ _00936_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_39_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout306 net181 net306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09811_ _01468_ _04490_ _04491_ _02598_ _04480_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_61_1388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09742_ _04380_ _04393_ _03182_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06954_ _01859_ _01867_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_138_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05905_ _00910_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09673_ _04358_ _02716_ _02766_ _03858_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10133__A1 _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06885_ _01716_ _01801_ _01802_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08877__A2 _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08624_ as2650.stack\[0\]\[3\] _03292_ _03293_ as2650.stack\[1\]\[3\] _03252_ _03326_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_96_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05836_ _00789_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_90_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_316 io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_77_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_327 la_data_out[48] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_77_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_as2650_338 la_data_out[49] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_132_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08555_ as2650.stack\[11\]\[1\] _03244_ _03246_ as2650.stack\[10\]\[1\] _03259_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_05767_ _00773_ _00777_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_166_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08629__A2 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07506_ _02315_ net370 _02309_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07837__B1 _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _01297_ _01702_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05698_ _00709_ _00710_ _00711_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10987__A3 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07437_ net281 _02256_ _02249_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11071__I _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07368_ _02191_ _02204_ _02205_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09107_ _03702_ _03796_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06319_ _01240_ _01246_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_116_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07299_ net293 _02137_ _02128_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_108_1521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06812__A1 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08380__I _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ _02474_ _03729_ _01367_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_148_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output174_I net174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_107_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11000_ _03817_ as2650.regs\[4\]\[6\] _05428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07907__A4 _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10372__A1 _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09109__A3 _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07724__I _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08317__B2 net211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_102_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08868__A2 _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06879__A1 _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10150__I _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_116_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09817__A1 _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_1546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11764_ _00543_ clknet_leaf_6_wb_clk_i as2650.stack\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_161_Right_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_81_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10715_ as2650.stack\[8\]\[3\] _05191_ _05195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11695_ _00479_ clknet_leaf_96_wb_clk_i as2650.regs\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10646_ _04768_ _05146_ _05149_ _04785_ _05151_ _05152_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_0_153_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_133_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xrebuffer5 net352 net349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_94_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_7__leaf_wb_clk_i clknet_leaf_51_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10577_ _01939_ _05104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_125_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06803__A1 _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_1698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11129_ as2650.stack\[14\]\[13\] _05515_ _05517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_34_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08859__A2 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06670_ _01598_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_1468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05621_ _00626_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_91_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09808__A1 net214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08340_ _00634_ _03060_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_43_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08271_ _01506_ _01308_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_1393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07222_ _02073_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07153_ _02029_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06104_ _01050_ net240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07809__I _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08795__B2 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07084_ _01835_ _01980_ _01983_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06035_ _00767_ net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_144_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ _01450_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_09725_ _01564_ _03736_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06937_ _01841_ _01851_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__11066__I _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _04340_ _04341_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__A3 _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06868_ _01785_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_1823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_1557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08607_ _03301_ _03304_ _03307_ _03309_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_52_1811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05819_ _00814_ _00817_ net198 _00827_ _00734_ _00704_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_09587_ _03658_ _03741_ _04258_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06799_ _01719_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08538_ _01274_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08469_ _00831_ _03171_ _03178_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10500_ as2650.stack\[1\]\[3\] _05048_ _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output291_I net291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11480_ _00264_ clknet_leaf_50_wb_clk_i as2650.irqs_latch\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07038__A1 _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10431_ _01380_ _04865_ _05002_ _04864_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_85_1653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08786__A1 _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07719__I _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10362_ _04162_ _04782_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10293_ _04863_ _04868_ _04869_ _04727_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_131_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10345__A1 _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_1562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07210__A1 net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07454__I _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05772__B2 _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_122_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_122_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_83_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08710__B2 as2650.stack\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05702__I as2650.debug_psl\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11747_ _00000_ clknet_leaf_87_wb_clk_i as2650.chirpchar\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_1428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11678_ _00462_ clknet_leaf_24_wb_clk_i as2650.stack\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09018__A2 _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_133_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_1727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10629_ _05108_ _05135_ _05138_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_12_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08777__A1 _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10336__A1 _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07840_ _02606_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_32_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_142_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07771_ _01965_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09510_ _04194_ _01768_ _01747_ _04195_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06722_ _01637_ _01627_ _01646_ _01647_ net186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_56_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__A1 _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _04108_ _04126_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_4_4__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06653_ _01588_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05604_ as2650.indirect_target\[6\] _00599_ _00615_ as2650.PC\[6\] _00618_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_59_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09372_ _04047_ _04053_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06584_ as2650.cycle\[2\] _01532_ _01514_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_133_1477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09257__A2 _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08323_ _03006_ _01315_ _01299_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11064__A2 _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_1604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_151_Left_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08254_ _02974_ _02986_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10811__A2 _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ net102 _02060_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_127_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08185_ _02926_ _02928_ _02925_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07136_ _02014_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_82_1837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07067_ _01971_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_101_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput240 net240 requested_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input50_I ram_bus_in[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput251 net251 requested_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_101_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput262 net262 rom_bus_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06018_ _00793_ net192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_80_1561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput273 net273 wbs_dat_o[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput284 net284 wbs_dat_o[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput295 net295 wbs_dat_o[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XPHY_EDGE_ROW_160_Left_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10878__A2 _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__I _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_162_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output137_I net137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07969_ _02614_ _01764_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09708_ _04392_ _04393_ _01477_ _01529_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_78_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10980_ _05313_ _05412_ _05405_ as2650.regs\[0\]\[1\] _05413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09639_ _02801_ _04322_ _04324_ _02626_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_97_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11601_ _00385_ clknet_leaf_88_wb_clk_i as2650.stack\[2\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10263__B1 _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11532_ _00316_ clknet_leaf_0_wb_clk_i as2650.stack\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11463_ _00247_ clknet_leaf_44_wb_clk_i as2650.PC\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_115_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_1401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08759__A1 _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10414_ _03120_ _04934_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_85_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11394_ _00178_ clknet_leaf_123_wb_clk_i as2650.chirp_ptr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10345_ _04815_ _04919_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_72_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _04803_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09184__A1 _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_124_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08931__A1 _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06388__I3 _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_124_wb_clk_i_I clknet_4_3__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_100_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_20_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07670__A1 net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07422__A1 net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09990_ _04595_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_110_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08941_ as2650.debug_psl\[0\] as2650.debug_psl\[3\] _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10513__I _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08872_ as2650.stack\[7\]\[12\] _03495_ _03514_ as2650.stack\[6\]\[12\] _03565_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07823_ _01092_ _02577_ _02589_ _02591_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_58_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07754_ _02486_ _02507_ _02514_ _02522_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09478__A2 _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06705_ _01631_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_17_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06866__C _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07685_ _02449_ _02457_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_79_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08150__A2 _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09424_ _00764_ _00774_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06438__I _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06636_ _01572_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_94_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08854__S _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09355_ _04039_ _04040_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06567_ as2650.ext_io_addr\[6\] _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_48_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08306_ _02998_ _02937_ _03030_ _03010_ _03031_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_35_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09286_ _03967_ _03971_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06498_ _01262_ _01459_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_1_1645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09650__A2 _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08237_ _02968_ _02970_ _02971_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06464__A2 _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ as2650.instruction_args_latch\[13\] _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_43_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09402__A2 _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10548__A1 _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_108_wb_clk_i clknet_4_8__leaf_wb_clk_i clknet_leaf_108_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07119_ net105 _02006_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06216__A2 _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08610__B1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08099_ as2650.ivectors_base\[5\] _02744_ _02850_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10130_ _01083_ _01573_ _03742_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_101_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output254_I net254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_164_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05975__A1 _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09166__A1 _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10061_ _01946_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09705__A3 _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08913__A1 _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10720__A1 _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10963_ _05396_ _05397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_104_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_104_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08141__A2 _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10894_ _05315_ _04902_ _05332_ _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08563__I _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08444__A3 _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11515_ _00299_ clknet_leaf_53_wb_clk_i net142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_81_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_74_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11446_ _00230_ clknet_leaf_38_wb_clk_i as2650.ivectors_base\[6\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10539__A1 _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11377_ _00173_ clknet_leaf_63_wb_clk_i as2650.insin\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07955__A2 _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06811__I _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10328_ _04881_ _04843_ _04903_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05966__A1 _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ _01747_ _04774_ _04836_ _04779_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__08939__S _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07707__A2 _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08904__A1 _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_1_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07642__I _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09704__I0 net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07470_ _02073_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06143__A1 _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06421_ _01346_ _01377_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_147_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06694__A2 _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11019__A2 _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _03825_ _03632_ _03826_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06352_ _01138_ _01301_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_6_wb_clk_i vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_56_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10778__A1 _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06283_ _01254_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07643__A1 net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ _03701_ _03705_ _03760_ _03761_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_72_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07089__I _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08022_ _02000_ _02777_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08199__A2 _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07817__I _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09973_ _01737_ _04596_ _04599_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_1427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08924_ _03613_ _03615_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_110_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08855_ _01920_ _03351_ _03548_ _03312_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07806_ net139 _01157_ _02574_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__08371__A2 _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ _01893_ _03347_ _03193_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_169_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05998_ _00969_ _00998_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_19_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input13_I bus_in_serial_ports[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07737_ _02505_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08659__B1 _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_157_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07668_ wb_counter\[29\] wb_counter\[30\] _02440_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_165_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_157_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09407_ _03916_ _03924_ _04092_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06619_ wb_debug_cc _01560_ _01540_ _01562_ _01556_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07599_ wb_counter\[16\] _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_153_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09338_ _04020_ _04022_ _04023_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08383__I _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06437__A2 _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_1464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09269_ _03944_ _03953_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08831__B1 _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11300_ _00096_ clknet_leaf_143_wb_clk_i net297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11231_ _00027_ clknet_leaf_133_wb_clk_i as2650.stack\[12\]\[10\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11194__A1 _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11162_ as2650.stack\[13\]\[9\] _05536_ _05538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06631__I _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10941__A1 _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10113_ _04663_ _04687_ _04692_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11093_ _05493_ _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_101_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10044_ _04626_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xhold50 net102 net394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_14__leaf_wb_clk_i clknet_leaf_76_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_106_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold61 net434 net405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold72 net459 net416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold83 _02005_ net427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_67_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold94 wbs_dat_i[11] net440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10946_ _04210_ _05303_ _05380_ _05381_ _05382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_133_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10877_ _05315_ _04872_ _05316_ _05317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08293__I as2650.instruction_args_latch\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06806__I _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11429_ _00213_ clknet_leaf_52_wb_clk_i as2650.instruction_args_latch\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07928__A2 _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08050__A1 _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10393__C1 _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11159__I _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06970_ _01882_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_52_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09852__I _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input5_I bus_in_gpios[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05921_ _00613_ _00616_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09550__A1 _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08353__A2 _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08640_ _02733_ _03064_ _03228_ _03341_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_05852_ as2650.regs\[3\]\[1\] _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06364__A1 _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10160__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _01762_ _02482_ _03241_ _03274_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05783_ _00793_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_89_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09302__A1 _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07522_ _02327_ _02328_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_147_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10999__A1 _05369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09853__A2 _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07453_ _02081_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06404_ net206 _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07321__B _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07384_ _02191_ _02217_ _02219_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09123_ _03755_ _03362_ _03723_ net215 _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06335_ _01243_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_33_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_1426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09054_ _03741_ _03742_ _03743_ _03745_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_142_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06266_ _01237_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_108_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08005_ _02712_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_1747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07219__I1 net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_635 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06197_ _01115_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08041__A1 _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__A2 _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09956_ _01629_ _04588_ _03051_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08907_ _02575_ _03589_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09887_ _04525_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_77_1533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08838_ _02762_ _03509_ _03532_ _03278_ _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10151__A2 _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output217_I net217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08769_ _03210_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_90_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10800_ _05100_ _05243_ _05247_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_155_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11780_ _00559_ clknet_leaf_4_wb_clk_i as2650.stack\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07155__I0 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10731_ as2650.stack\[8\]\[9\] _05203_ _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10662_ as2650.regs\[1\]\[7\] _05162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06626__I _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_123_wb_clk_i clknet_4_9__leaf_wb_clk_i clknet_leaf_123_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07607__A1 net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10148__I _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10593_ _05115_ _05116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11167__A1 _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07457__I _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06361__I _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11214_ _05469_ _05568_ _05570_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_92_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10914__A1 net191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08583__A2 _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09780__A1 _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11145_ _05445_ _05522_ _05527_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06594__A1 _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09672__I _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__05906__S _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11076_ as2650.regs\[7\]\[1\] _05484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08335__A2 _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _04633_ _04625_ _04634_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10142__A2 _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08099__A1 as2650.ivectors_base\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_13__f_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07146__I0 net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10929_ _04964_ _05364_ _05365_ _05276_ _05366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_168_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_99_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09599__A1 _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10058__I _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06120_ _01090_ _01091_ _01092_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__08271__A1 _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06051_ _01034_ net256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_129_1493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08023__A1 as2650.indirect_target\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08023__B2 _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__A1 _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09810_ _02560_ _04479_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_39_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08399__S _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10381__A2 _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09741_ _04425_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_06953_ _01787_ _01865_ _01866_ _01798_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09523__A1 _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05904_ _00708_ _00908_ _00909_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09672_ _01349_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_94_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06884_ as2650.stack\[12\]\[3\] _01739_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10133__A2 _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08623_ as2650.stack\[3\]\[3\] _03264_ _03254_ as2650.stack\[2\]\[3\] _03325_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05835_ _00692_ _00842_ _00843_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_94_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_317 irq[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_328 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_08554_ _03247_ _03253_ _03255_ _03257_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07137__I0 net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05766_ _00705_ _00774_ _00776_ _00736_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xwrapped_as2650_339 la_data_out[50] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07505_ net101 _02307_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07837__B2 _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08485_ _00597_ _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05697_ _00709_ as2650.regs\[6\]\[7\] _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_1835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07436_ _02244_ wb_counter\[23\] _02263_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07367_ net270 _02197_ _02188_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _03705_ _03795_ _03785_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06318_ _01248_ _01273_ _01288_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_60_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08262__A1 _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08262__B2 net203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07298_ _02114_ wb_counter\[5\] _02143_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_1819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09037_ _03587_ _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06249_ _01221_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_130_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_148_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08565__A2 _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09939_ _04571_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08317__A2 _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08868__A3 _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07128__I0 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07740__I _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11763_ _00542_ clknet_leaf_5_wb_clk_i as2650.stack\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ _05080_ _05189_ _05194_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_81_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11694_ _00478_ clknet_leaf_96_wb_clk_i as2650.regs\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_137_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10645_ as2650.regs\[1\]\[0\] _05152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_133_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer6 net349 net350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10576_ _05102_ _05095_ _05103_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_94_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06803__A2 _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_90_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_91_wb_clk_i clknet_4_10__leaf_wb_clk_i clknet_leaf_91_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08556__A2 _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09753__A1 _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_20_wb_clk_i clknet_4_1__leaf_wb_clk_i clknet_leaf_20_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07915__I _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11128_ _05469_ _05514_ _05516_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_34_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06319__A1 _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ _05469_ _05470_ _05472_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_88_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10115__A2 _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_4_6__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05620_ as2650.page_reg\[0\] _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_8_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07819__A1 _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08270_ _01265_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_28_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07221_ net66 _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_89_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_rebuffer3_I _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold110_I wbs_dat_i[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07152_ net74 net124 _02025_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06103_ _01055_ net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__08414__C _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__A1 as2650.stack\[4\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07083_ as2650.stack\[11\]\[5\] _01981_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_1710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06034_ _00730_ net218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06270__A3 _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_143_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07755__B1 _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08430__B _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07985_ as2650.indirect_target\[3\] _02723_ _02738_ _02742_ _02743_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_96_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09724_ _04270_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06936_ _01843_ _01847_ _01850_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_39_1612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10106__A2 _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09655_ _02726_ _01643_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_1525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06867_ _01722_ _01723_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_97_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ as2650.stack\[15\]\[2\] _03308_ _03142_ as2650.stack\[14\]\[2\] _03298_ _03309_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05818_ _00826_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_132_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09586_ _04255_ _04256_ _04271_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06798_ as2650.PC\[0\] _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_136_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08537_ _03224_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10409__A3 _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05749_ _00694_ _00759_ _00760_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11082__I _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08483__A1 _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07286__A2 _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ as2650.ivectors_base\[7\] _03172_ _03175_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10290__A1 _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07419_ net278 _02225_ _02249_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08399_ _03113_ _03119_ _02552_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10430_ _02913_ _01363_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06904__I _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07038__A2 _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08235__B2 net198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output284_I net284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08786__A2 _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10361_ _01804_ _04932_ _04935_ _04876_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_104_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_1390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06261__A3 _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10292_ _01410_ _04758_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_1362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09735__A1 _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07735__I _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_70_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__05772__A2 _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_122_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06721__A1 net249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07470__I _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_114_wb_clk_i_I clknet_4_10__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07277__A2 _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11746_ _00530_ clknet_leaf_115_wb_clk_i as2650.stack\[0\]\[15\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09671__B1 _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11677_ _00461_ clknet_leaf_18_wb_clk_i as2650.stack\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10628_ as2650.stack\[7\]\[13\] _05136_ _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07029__A2 _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_1430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10559_ _05090_ _05085_ _05091_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10584__A2 _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_1514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07770_ _02509_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_153_wb_clk_i_I clknet_4_0__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06721_ net249 _01617_ _01600_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09440_ _04090_ _04091_ _04107_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_56_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06652_ _01239_ _01587_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_91_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05603_ as2650.indirect_target\[5\] _00598_ _00614_ as2650.PC\[5\] _00617_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_8_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09371_ _04025_ _04043_ _04056_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06583_ _01529_ _01273_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_75_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08322_ _03000_ _02992_ _03002_ net212 _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_150_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08465__A1 _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08253_ as2650.instruction_args_latch\[5\] _02975_ _02985_ _02981_ _02986_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_89_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07204_ _02058_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08184_ _02927_ _02917_ _02922_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10024__A1 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__A1 net227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ _02019_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08768__A2 _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06779__A1 _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07066_ _01961_ _01962_ _01970_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput230 net230 last_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_144_1574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07440__A2 wb_counter\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput241 net241 requested_addr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput252 net252 requested_addr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_1513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06017_ _00758_ net193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_100_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput263 net263 rom_bus_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_140_1449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput274 net274 wbs_dat_o[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput285 net285 wbs_dat_o[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input43_I irqs[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput296 net296 wbs_dat_o[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_162_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07968_ _02725_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_138_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09707_ net8 net16 net32 net24 as2650.ext_io_addr\[7\] _04384_ _04393_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_06919_ _01834_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07899_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_97_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08386__I _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09638_ _01806_ _02465_ _04323_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07290__I _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09569_ _01031_ _01388_ _01501_ _01390_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_112_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11600_ _00384_ clknet_leaf_122_wb_clk_i as2650.stack\[2\]\[14\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09653__B1 _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11531_ _00315_ clknet_leaf_0_wb_clk_i as2650.stack\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_22_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11462_ _00246_ clknet_leaf_44_wb_clk_i as2650.PC\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06634__I _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_115_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10413_ _04364_ _04843_ _04985_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_145_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11393_ _00177_ clknet_leaf_36_wb_clk_i as2650.cpu_hidden_rom_enable vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10344_ _01397_ _04917_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_72_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09708__A1 _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10275_ _04733_ _04850_ _04851_ _04740_ _01769_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_128_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08070__B _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_1807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11729_ _00513_ clknet_leaf_83_wb_clk_i as2650.regs\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06473__A3 _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07670__A2 _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09947__A1 _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__A2 _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08940_ _03628_ _03630_ _03631_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_102_1709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07375__I _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08871_ as2650.stack\[0\]\[12\] _03516_ _03517_ as2650.stack\[1\]\[12\] _02505_ _03564_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_97_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07822_ _02590_ _02576_ _02567_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_93_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07753_ as2650.stack\[4\]\[13\] _02493_ _02500_ as2650.stack\[5\]\[13\] _02521_ _02522_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_75_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06704_ _01605_ _01371_ _01630_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_07684_ net231 _01638_ _01654_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_1517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09423_ _04099_ _04102_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_1539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06635_ _01098_ _00968_ _00997_ _01074_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_165_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09354_ _04020_ _04022_ _04030_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_06566_ _01518_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_136_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08438__A1 _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10245__A1 _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08305_ _03021_ _02627_ _03022_ net208 _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09285_ _03969_ _03970_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07110__A1 _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06497_ _01266_ _01191_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_133_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08236_ as2650.instruction_args_latch\[3\] _02955_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05672__A1 _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08167_ _02911_ _02912_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10548__A2 _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07118_ wb_feedback_delay _02005_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ _02837_ _02845_ _02847_ _02849_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08610__A1 _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07049_ _01930_ _01954_ _01955_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_164_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_148_wb_clk_i clknet_4_2__leaf_wb_clk_i clknet_leaf_148_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10060_ _04655_ _04656_ _04658_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_1399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output247_I net247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09705__A4 _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_10_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_1387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06924__A1 _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_3_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10962_ _05147_ _05395_ _03816_ _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_74_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08677__B2 as2650.stack\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10893_ _04881_ _05315_ _05332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06152__A2 _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08429__A1 _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10236__A1 _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11514_ _00298_ clknet_leaf_53_wb_clk_i net141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_78_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08444__A4 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05663__A1 _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11445_ _00229_ clknet_leaf_38_wb_clk_i as2650.ivectors_base\[5\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_123_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10539__A2 _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11376_ _00172_ clknet_leaf_63_wb_clk_i as2650.insin\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_156_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10614__I _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10327_ _04844_ _04902_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05708__I _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _03498_ _04775_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08904__A2 _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10189_ _04767_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__05718__A2 _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07923__I _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10711__A2 _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09704__I1 net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08668__A1 _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06539__I _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06420_ _01383_ _01360_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10227__A1 _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06351_ _01268_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11180__I _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09070_ _00732_ _02677_ _03708_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06282_ _01253_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_115_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08021_ _02638_ _02774_ _02776_ _02705_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09396__A2 _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09972_ as2650.stack\[4\]\[0\] _04598_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05957__A2 _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09148__A2 _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08923_ _00833_ _03586_ _03614_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08854_ _03542_ _03547_ _02551_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07805_ net63 net139 _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08785_ _03235_ _03454_ _03481_ _03234_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_05997_ _00997_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_135_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07736_ _02504_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_7_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07667_ _02332_ _02444_ _02445_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_157_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_157_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06618_ as2650.insin\[6\] _01561_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09406_ _03919_ _03923_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07598_ _02357_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06549_ _01503_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09337_ _04018_ _04019_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_1787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09268_ _03953_ _03944_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output197_I net197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08219_ _02904_ _02953_ _02956_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_112_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09199_ _03874_ _03883_ _03884_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_69_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11230_ _00026_ clknet_leaf_133_wb_clk_i as2650.stack\[12\]\[9\] vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07398__A1 net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11161_ _05459_ _05535_ _05537_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10112_ as2650.stack\[3\]\[15\] _04688_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09139__A2 _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11092_ _01685_ _05186_ _04622_ _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_105_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10043_ _04624_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_101_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_1815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08839__I _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08898__A1 _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold40 net444 net384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__07743__I _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xhold51 net455 net395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold62 net460 net406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_106_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold73 net443 net417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold84 wbs_we_i net428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_TAPCELL_ROW_67_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold95 wbs_dat_i[12] net441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_TAPCELL_ROW_67_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_1534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10945_ _04169_ _04781_ _05341_ _05381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_5__leaf_wb_clk_i clknet_leaf_45_wb_clk_i vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_hold99_I wbs_dat_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_1608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _04842_ _04844_ _05316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_1843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05884__A1 _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__A1 _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07918__I _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11428_ _00212_ clknet_leaf_55_wb_clk_i as2650.instruction_args_latch\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_65_1663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06822__I _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11185__A2 _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11359_ _00155_ clknet_leaf_102_wb_clk_i wb_counter\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10393__B1 _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05920_ _00660_ _00924_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_52_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05851_ _00588_ _00658_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06269__I _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08570_ _03242_ _03273_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05782_ _00792_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_72_1623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07521_ _02091_ _02101_ _02108_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_1679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09302__A2 _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07313__A1 net182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07452_ _02190_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05875__A1 _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06403_ _00886_ net206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_169_1422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07383_ net272 _02197_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09066__A1 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09122_ _03806_ _03810_ _03051_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06334_ _01249_ _01302_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_112_1690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08813__A1 _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09053_ _03744_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_06265_ _01236_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_72_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08004_ _02572_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07828__I _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06732__I _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06196_ _01168_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_13_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07919__A3 _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08041__A2 _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09955_ net222 _04586_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08906_ _01346_ _01227_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09886_ _01928_ _04539_ _04544_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08837_ _01469_ _03511_ _03531_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_1822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_159_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ as2650.stack\[0\]\[8\] _03261_ _03262_ as2650.stack\[1\]\[8\] _03464_ _03465_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_TAPCELL_ROW_101_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output112_I net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07719_ _02487_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08699_ _01846_ _03347_ _03372_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07155__I1 net125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11100__A2 _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10730_ _05094_ _05202_ _05204_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06907__I _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10661_ _04986_ _05156_ _05157_ _04989_ _05158_ _05161_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09057__A1 net188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10592_ _05114_ _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08804__A1 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__A1 _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11213_ as2650.stack\[9\]\[12\] _05569_ _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_1403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11144_ as2650.stack\[13\]\[2\] _05524_ _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06594__A2 _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11075_ _05163_ _05480_ _05482_ _05483_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_95_1601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_hold14_I net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ as2650.stack\[10\]\[3\] _04627_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08335__A3 _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_4_1__leaf_wb_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08740__B1 _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08099__A2 _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09296__A1 _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07146__I1 net136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10928_ _04171_ _04778_ _05365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__05721__I net345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05857__A1 _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09048__A1 _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10859_ as2650.regs\[4\]\[1\] _05288_ _05300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_99_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06050_ net66 _01033_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_2_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08559__B1 _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09740_ _02813_ _04372_ _04380_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06952_ _01860_ _01793_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends

