* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i wb_rst_i
XFILLER_100_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7406__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__I0 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7963_ _1644_ _3316_ _3274_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _1613_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7894_ _1564_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8657__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6845_ _2244_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8382__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _0407_ _2188_ _2193_ as2650.r123_2\[1\]\[2\] _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8515_ _3789_ _3804_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5727_ _1260_ _1073_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7256__I _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__A2 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6160__I _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8446_ as2650.r123\[2\]\[3\] _3741_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5658_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7893__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ _4189_ _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8377_ _1240_ _1295_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7893__B2 _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _1115_ _1134_ _1136_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7328_ _2700_ _2702_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7645__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6448__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7259_ _1581_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__A1 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6999__A3 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__S _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8070__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5959__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6335__I _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6923__A3 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8125__A2 _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6070__I _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7636__A1 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7939__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8061__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ as2650.holding_reg\[4\] _4166_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_92_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4891_ _0382_ _0429_ _0449_ _4059_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7167__A3 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8364__A2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _2078_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8460__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6375__A1 _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6561_ _2012_ _2013_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_125_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7076__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8116__A2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8300_ _0876_ _3189_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5512_ _0890_ _0908_ _0909_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6492_ _1771_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8231_ _3526_ _2808_ _3527_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5443_ _0940_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8162_ _3470_ _3475_ _3155_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5350__A2 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ as2650.stack\[2\]\[8\] _0920_ _0927_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7627__A1 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7113_ _1085_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4325_ _3901_ _3905_ _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8093_ _2632_ _2734_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7044_ _0320_ _2422_ _2435_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__A2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7946_ _1564_ _1356_ _3299_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7877_ _3158_ _1345_ _3235_ _1550_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _1409_ _1267_ _2220_ _2236_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6759_ as2650.r123_2\[0\]\[6\] _2154_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4403__I as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__A4 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6118__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8429_ _3731_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__A1 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8822__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8043__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__I _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5409__I _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6109__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7624__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6124__A4 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5332__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__A1 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7609__B2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__A1 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5090_ _0378_ _4230_ _0369_ _0542_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_111_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4983__I _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6832__A2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8034__A1 as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8585__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7800_ _1585_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8780_ _0179_ clknet_3_3_0_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5992_ _1216_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7731_ _2621_ _3073_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7662_ _1188_ _2943_ _2914_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6348__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4874_ _4014_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8123__C _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _1360_ _1812_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6899__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ _1177_ _2914_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6544_ _0454_ _1900_ _1857_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7962__C _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7848__A1 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6475_ _0665_ _0614_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8214_ _2757_ _2824_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5426_ _0957_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6520__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8845__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4531__B1 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8145_ _3434_ _3457_ _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5357_ _0894_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4308_ _3888_ _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8273__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8076_ _3191_ _4062_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5288_ _0753_ _0675_ _0752_ _0756_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5087__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7027_ _2420_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6823__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8025__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7929_ _0574_ _3161_ _3163_ _2891_ _1563_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_70_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5229__I _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5562__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7839__A1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8264__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__I _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8016__A1 as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4308__I _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8319__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8718__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7782__C _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8868__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4590_ _3946_ _4170_ _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7354__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6502__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5305__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _4281_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6191_ _1644_ _1685_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8255__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5142_ _0699_ _0700_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_97_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6266__B1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _0631_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__I _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4816__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8007__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7022__C _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8832_ _0231_ clknet_leaf_20_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8763_ _0162_ clknet_leaf_0_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5975_ _1192_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7714_ _1396_ _3077_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4926_ _4172_ _0472_ _0487_ _4148_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8694_ _0093_ clknet_leaf_24_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7645_ _1190_ _2608_ _3012_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4857_ _0417_ _3895_ _4103_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8191__B1 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7576_ _2613_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4788_ net7 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6741__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6527_ _1934_ _1938_ _1980_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7297__A2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8494__A1 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6458_ as2650.r123_2\[2\]\[1\] _1830_ _1913_ _1862_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5409_ _0310_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6389_ _4206_ _1813_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8128_ _2483_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8246__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7049__A2 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8309__B _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8059_ _2136_ _3327_ _3376_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5480__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7221__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6024__A3 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4572__B _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A1 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8237__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7123__B _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__I _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7460__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7349__I _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6253__I _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _1282_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5774__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7793__B _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4711_ _4016_ _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5691_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7430_ _2766_ _2787_ _2799_ _2800_ _2802_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_72_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4642_ _4222_ _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5526__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8401__C _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _4268_ _4082_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4573_ _4143_ _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _4197_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7279__A2 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7292_ _2666_ _2629_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8228__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _1666_ _4270_ _0656_ _1667_ _1537_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_69_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ _0456_ _0654_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__A4 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5056_ _0609_ _0610_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7968__B _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__A1 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8815_ _0214_ clknet_leaf_33_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7203__A2 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7259__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8746_ _0145_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5958_ as2650.stack\[1\]\[8\] _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4909_ _4189_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5889_ _1245_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8677_ _0076_ clknet_leaf_47_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7628_ _1189_ _2995_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5517__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6714__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7559_ _2925_ _2880_ _2927_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6190__A2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7878__B _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6953__A1 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A2 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6181__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__I _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8458__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A1 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7681__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A2 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__A3 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5444__B2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8463__I _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6930_ _1575_ _1373_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7197__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6861_ _2063_ _2248_ _2264_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8600_ _2492_ _3881_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5812_ _1326_ _1342_ _1343_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6792_ _2208_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5743_ _1272_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8531_ _0349_ _0478_ _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5674_ as2650.pc\[11\] _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8462_ _2459_ _1727_ _3755_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7413_ _2777_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _4203_ _3964_ _4205_ _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8393_ _3080_ _3697_ _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7344_ _2715_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4556_ _4134_ _4135_ _4136_ _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_132_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7275_ _0976_ _2650_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4487_ net5 _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _1148_ _1704_ _1708_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6157_ net1 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _0667_ _3895_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7698__B _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _1580_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _4211_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7188__A1 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6935__A1 _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8729_ _0128_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 net20 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput31 net31 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7452__I _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput42 net42 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7663__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7401__B _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7274__S1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7351__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A2 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4410_ _3940_ _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5390_ _0943_ as2650.stack\[5\]\[8\] as2650.stack\[4\]\[8\] _0946_ _0947_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_67_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _3917_ _3921_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7103__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7060_ _1167_ _2433_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7654__A2 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _0532_ _0754_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7406__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__I1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7962_ _1561_ _1361_ _3313_ _3315_ _1684_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5610__I _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5968__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6090__A1 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6913_ _2226_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7893_ _1210_ _3161_ _3163_ _2799_ _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_78_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ as2650.addr_buff\[1\] _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6917__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7965__C _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6775_ _1965_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8514_ _1841_ _2992_ _2375_ _3756_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5726_ _3901_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8445_ _3738_ _1989_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7342__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5657_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6145__A2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4608_ _4188_ _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8376_ _3044_ _3681_ _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5588_ as2650.stack\[5\]\[1\] _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4539_ _3958_ _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7327_ as2650.stack\[2\]\[1\] _0919_ _0927_ _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7272__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7645__A2 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4459__A2 _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ as2650.stack\[0\]\[4\] _1696_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7189_ _2562_ _2563_ _2567_ _2455_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5408__A1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7221__B _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8070__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5959__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8601__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6908__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8751__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__I _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7333__A1 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4698__A2 _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8278__I _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4942__I0 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7636__A2 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7910__I as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8597__B1 _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6072__A1 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _0450_ _0451_ _0381_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7572__A1 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6375__A2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6261__I _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _4097_ _0574_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5511_ _4197_ _0904_ _1060_ _0894_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6491_ _1916_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8230_ _2408_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5442_ _0943_ as2650.stack\[5\]\[10\] as2650.stack\[4\]\[10\] _0946_ _0997_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8161_ _3402_ _3472_ _3474_ _3443_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5373_ as2650.stack\[1\]\[8\] as2650.stack\[0\]\[8\] _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5605__I _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4324_ _3904_ _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8092_ _3407_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7043_ _1600_ _2419_ _2432_ _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_86_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8624__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8052__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7945_ _1233_ _3161_ _3163_ _2939_ _3159_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_83_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7876_ _3160_ _4092_ _3234_ _1567_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6827_ _1286_ _2235_ _3985_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7563__A1 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7563__B2 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5709_ _3943_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7315__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6118__A2 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6689_ _1163_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8428_ _4034_ _1397_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8359_ _3402_ _3665_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7079__B1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7618__A2 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5629__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8291__A2 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8043__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4604__A2 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A2 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7857__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6030__B _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__A2 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6832__A3 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8797__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6256__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8034__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__A3 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5991_ _1490_ _1483_ _1491_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ _3070_ _3073_ _3093_ _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4942_ as2650.r123\[0\]\[3\] as2650.r123_2\[0\]\[3\] _3887_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7661_ _1196_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7545__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6348__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4873_ _0427_ _0354_ _0355_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4504__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6612_ _2063_ _1847_ _1848_ _0662_ _1850_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_123_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6899__A3 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7592_ _1544_ _2876_ _2958_ _2960_ _2733_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_6543_ _1839_ _1994_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7848__A2 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _1927_ _1928_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8213_ _3519_ _3524_ _1314_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5425_ _0970_ _0974_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5335__I _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6520__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4531__A1 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5356_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8144_ _4269_ _4232_ _4235_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4531__B2 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4307_ _3887_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8075_ _1314_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8273__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5087__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7026_ _1600_ _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ as2650.psu\[5\] _3210_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7536__A1 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _2251_ _1643_ _1577_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4414__I _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7839__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6511__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8264__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_39_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6275__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7472__B1 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A3 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8016__A2 _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7775__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4324__I _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8878__D _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0626_ _0752_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6190_ _1561_ _1360_ _1683_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5141_ _0365_ _0401_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8255__A2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__B2 _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _0532_ _0533_ _0527_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__A2 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__B _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8831_ _0230_ clknet_leaf_28_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8415__B _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7766__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7766__B2 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8762_ _0161_ clknet_leaf_78_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _1237_ _1473_ _1477_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7713_ as2650.addr_buff\[3\] _3076_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4925_ _0473_ _0475_ _0481_ _0331_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7518__A1 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8693_ _0092_ clknet_leaf_74_wb_clk_i as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7644_ _2982_ _3008_ _3010_ _2991_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4856_ as2650.r123\[1\]\[4\] as2650.r123\[0\]\[4\] as2650.r123_2\[1\]\[4\] as2650.r123_2\[0\]\[4\]
+ _3882_ _3888_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8812__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8191__B2 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7575_ _2943_ _2897_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4787_ _0295_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__C _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4752__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ _0667_ _0615_ _1939_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _1899_ _1912_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5408_ as2650.r123\[0\]\[1\] _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6388_ _1823_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ _3423_ _3424_ _3440_ _3441_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7280__I _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _4192_ _4190_ _4193_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6257__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8058_ as2650.stack\[7\]\[6\] _3324_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _1288_ _2404_ _2291_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6009__A1 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__A1 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5232__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7455__I _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A2 _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5299__A2 _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7123__C _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__I _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7748__A1 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8835__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__A1 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _4284_ _4289_ _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ as2650.pc\[13\] _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4641_ _4221_ _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7360_ _1268_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4572_ _4148_ _4152_ _4146_ _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6311_ _3969_ _1071_ _4015_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7291_ _1429_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6242_ _1249_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8228__A2 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ as2650.psl\[6\] _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5613__I _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _4042_ _0679_ _0683_ _4277_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5055_ _4050_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7739__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__I _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8814_ _0213_ clknet_leaf_34_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5488__C _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6411__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8745_ _0144_ clknet_leaf_61_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4973__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8676_ _0075_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8164__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8164__B2 _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7627_ _2994_ _2914_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4839_ _4049_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6714__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7911__A1 _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4725__A1 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _2925_ _2880_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6509_ _0349_ _1950_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7489_ _2857_ _0560_ _2859_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8708__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7690__A3 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__I _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6650__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5398__C _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5756__A3 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7185__I _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7902__A1 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6705__A2 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8458__A2 _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6469__A1 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A2 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__B _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6529__I _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7969__A1 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__C _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6641__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _2263_ _2253_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5811_ net43 _1333_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ as2650.r123\[3\]\[0\] _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8530_ _0348_ _0478_ _3817_ _4289_ _3818_ _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5742_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8461_ _3754_ _1726_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5673_ _1126_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7412_ _2780_ _2782_ _2783_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4512__I _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4707__A1 _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4204_ _3956_ _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8392_ _3044_ _3681_ _3081_ _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7343_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__A2 _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ as2650.holding_reg\[0\] _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7274_ as2650.stack\[3\]\[0\] as2650.stack\[0\]\[0\] as2650.stack\[1\]\[0\] as2650.stack\[2\]\[0\]
+ _0915_ _0916_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4486_ _3954_ _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__B _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6225_ as2650.stack\[1\]\[3\] _1706_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6156_ as2650.psu\[3\] _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5107_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6087_ _1320_ _1390_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _0316_ _0548_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8385__A1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7188__A2 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6989_ _2343_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6902__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8728_ _0127_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8659_ _0058_ clknet_leaf_32_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__I _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__I _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput32 net32 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput43 net43 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6349__I _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8680__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4882__B1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6926__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6968__B _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6154__A3 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__I _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ as2650.addr_buff\[7\] _3920_ _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7103__A2 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8300__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6259__I _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5163__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6010_ _0522_ _0630_ _0845_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6614__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7961_ _2156_ _2976_ _3314_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6912_ _0878_ _2309_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7892_ _1651_ _3248_ _3249_ _0902_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6917__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4928__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6774_ _2190_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8119__A1 _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8513_ _1590_ _3802_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5725_ _1250_ _1253_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7039__B _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8444_ _0396_ _3733_ _3743_ _3744_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5656_ as2650.pc\[9\] _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _4165_ _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5353__A1 _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8375_ _3048_ _3680_ _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5587_ _1122_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7326_ as2650.stack\[1\]\[1\] as2650.stack\[0\]\[1\] _0928_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4538_ _3971_ _4118_ _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7257_ _1094_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ _4049_ _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _1148_ _1694_ _1698_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7188_ _2437_ _2369_ _2565_ _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _1631_ _1634_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4417__I _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6632__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8530__B2 _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5344__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4942__I1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7097__A1 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6079__I _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7412__B _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8597__A1 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8597__B2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8349__A1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__B _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5510_ _1059_ _0957_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ _1918_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4997__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5441_ as2650.stack\[2\]\[10\] _0920_ _0927_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8160_ _2717_ _3473_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5372_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _2494_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7088__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__B1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4323_ _3902_ _3903_ _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8091_ _2678_ _2337_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _1532_ _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__B1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8588__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7260__A1 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7944_ net27 _1388_ _3298_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7875_ _3213_ _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7548__I _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _3973_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6757_ _1048_ _0957_ _1054_ _2171_ _2153_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_91_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _1240_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _2130_ _2131_ _2132_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7315__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8512__A1 _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8427_ _3729_ _3730_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5326__A1 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _1150_ _1179_ _1180_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__I _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5877__A2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8358_ net50 _3664_ _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7079__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__B2 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7309_ net5 _4046_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8289_ net34 _3389_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5629__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8579__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7886__C _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6362__I _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8503__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6109__A3 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6817__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__A4 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ as2650.stack\[2\]\[10\] _1488_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7793__A2 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4941_ _0499_ _0500_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7660_ _2681_ _3026_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4872_ _4072_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ _1652_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5556__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7591_ _2829_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6542_ _0410_ _1995_ _1834_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_9_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8420__C _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5308__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6473_ _1883_ _1891_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5616__I _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8212_ _0561_ _3192_ _3523_ _3922_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5424_ _0977_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8143_ _4232_ _4235_ _4269_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5355_ _4191_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4306_ _3886_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8074_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5286_ as2650.holding_reg\[7\] _0737_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8741__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6284__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7025_ _1573_ _1616_ _1617_ _3951_ _2418_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_60_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5492__B1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7927_ _1667_ _3164_ _0903_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7278__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5300__B _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7858_ _1529_ _3217_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7536__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _2216_ _2217_ _1293_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7789_ _2460_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8497__B1 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6275__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7472__B2 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A4 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7897__B _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A1 _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7775__A2 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5786__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4605__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A2 _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__B1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6820__I _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8614__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7137__B _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5436__I _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8764__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ as2650.r0\[1\] _0612_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7463__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__A2 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5071_ _0519_ _0521_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5171__I _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8830_ _0229_ clknet_leaf_27_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7766__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8761_ _0160_ clknet_leaf_1_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ as2650.stack\[1\]\[14\] _1475_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7712_ as2650.addr_buff\[3\] _3076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4515__I as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _0482_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8692_ _0091_ clknet_leaf_74_wb_clk_i as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7643_ _2604_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7574_ as2650.pc\[7\] _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4786_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6525_ _1881_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4752__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6456_ _1833_ _1909_ _1911_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5701__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8126_ _2407_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5338_ _4200_ _0569_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_47_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7454__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6257__A2 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8057_ _2133_ _3327_ _3375_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ as2650.r0\[0\] _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _1303_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7206__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__I _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8637__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4440__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7509__A2 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8341__B _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8787__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5940__A1 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6248__A2 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__B1 as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7996__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6420__A2 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4431__A1 _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ _4220_ _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6184__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6184__B2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7920__A2 _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _4149_ _4150_ _4151_ as2650.holding_reg\[0\] _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5931__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _1500_ _1763_ _1767_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7290_ _1594_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _1715_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ as2650.psl\[5\] _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7436__A1 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _4042_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5998__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8426__B _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7739__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8813_ _0212_ clknet_leaf_28_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8744_ _0143_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5956_ _1463_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _0466_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8675_ _0074_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5887_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8164__A2 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7626_ _2943_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4838_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6175__A1 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7557_ _2926_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4769_ _4288_ _4294_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ _1950_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7488_ _2759_ _2858_ _2809_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7675__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _1870_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7291__I _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8109_ net52 _3400_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__A2 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7240__B _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__A2 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6402__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__A4 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7666__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__A2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7418__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_23_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8091__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8802__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8246__B _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4652__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8394__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5810_ _0993_ _1339_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6790_ _0843_ _2074_ _2207_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4404__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _1263_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8460_ _1535_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5672_ _0831_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7411_ _1087_ _2329_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _3957_ _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8391_ _3088_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7342_ as2650.pc\[2\] net7 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4554_ _4053_ _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__A1 _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7325__B _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7273_ _2648_ as2650.stack\[7\]\[0\] as2650.stack\[6\]\[0\] _0918_ _0953_ _2649_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4485_ _4065_ _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5624__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6224_ _1142_ _1704_ _1707_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7409__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _3885_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4891__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5106_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4891__B2 _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _4201_ _1581_ _1417_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _4282_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__A1 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6988_ _2159_ _1075_ _2381_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8727_ _0126_ clknet_leaf_26_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7286__I _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ as2650.stack\[0\]\[9\] _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8658_ _0057_ clknet_leaf_35_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__C _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6699__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _2665_ _2944_ _2976_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8589_ _1167_ _2436_ _3872_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput11 net11 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput22 net22 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput33 net33 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput44 net44 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5123__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8825__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4882__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A1 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5709__I _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6139__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__C _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7639__A1 _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__A2 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6311__A1 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8064__A1 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7811__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7960_ _2050_ _3162_ _3159_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4625__A1 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6911_ _2306_ _0733_ _2308_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_47_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7891_ _4095_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8367__A2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6842_ _4268_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_50_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8423__C _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6773_ _0313_ _2074_ _2196_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8119__A2 _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8512_ _3760_ _3801_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5724_ _1255_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7327__B1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7878__A1 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8443_ as2650.r123\[2\]\[2\] _3741_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5655_ _1187_ _1193_ _1195_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _4186_ _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8374_ _3018_ _3643_ _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8848__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5353__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7325_ as2650.stack\[3\]\[1\] _0934_ _0937_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4537_ _3974_ _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5354__I _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7256_ _4070_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6302__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _4048_ _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6207_ as2650.stack\[0\]\[3\] _1696_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7187_ _1298_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4399_ _3970_ _3975_ _3979_ _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6138_ as2650.psl\[6\] _1621_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _4110_ _0718_ _1361_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8070__A4 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8333__C _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4433__I _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7869__A1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8530__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7097__A2 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7412__C _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8597__A2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6095__I _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__I _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__C _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7021__A2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5032__A1 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8521__A2 _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5440_ as2650.stack\[1\]\[10\] as2650.stack\[0\]\[10\] _0929_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ _0915_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ _1687_ _1284_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8285__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7088__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4322_ net10 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_99_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8090_ _3405_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5099__A1 _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7041_ _2428_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6835__A2 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__A1 as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5902__I _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8037__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_1_1_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_opt_1_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8588__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7260__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7943_ _1668_ _3164_ _0903_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__I _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _0501_ _3162_ _0913_ _2751_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6825_ _4121_ _1304_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5349__I _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6756_ _2181_ _2182_ _2183_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_91_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8670__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _1093_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ as2650.stack\[4\]\[4\] _2124_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7315__A3 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8426_ net40 _3418_ _2402_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5638_ as2650.stack\[5\]\[7\] _1165_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5326__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8357_ _3636_ _3638_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5569_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7308_ _2678_ _1086_ _2680_ _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8276__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8276__B2 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8288_ _1168_ _3486_ _3597_ _3452_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7513__B _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7239_ _2612_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8579__A2 _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4428__I _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__A1 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6762__B2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5208__B _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6817__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6818__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__I _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8019__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4940_ _4256_ _4086_ _0306_ _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_92_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8693__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ _0429_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5169__I _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _0648_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7590_ _2956_ _2929_ _2957_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_92_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6753__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5556__A2 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7950__B1 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _1838_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7384__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _1886_ _1890_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6505__A1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5308__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ as2650.stack\[3\]\[9\] as2650.stack\[0\]\[9\] as2650.stack\[1\]\[9\] as2650.stack\[2\]\[9\]
+ _0929_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8211_ _2031_ _0594_ _3522_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_127_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8258__A1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8142_ _3978_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5354_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_142_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8258__B2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6269__B1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4305_ as2650.psl\[4\] _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8073_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6728__I _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5285_ _0809_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7024_ _3906_ _1612_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5492__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__C _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7926_ _3150_ _2062_ _3279_ _3280_ _3281_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_70_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _3158_ _4261_ _3215_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5079__I _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6808_ _1581_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6744__A1 _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7788_ _1234_ _2608_ _3149_ _3135_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _1555_ _0900_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7294__I _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5807__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__I _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8497__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8409_ _3485_ _3712_ _3713_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8249__A1 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5542__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7224__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8421__A1 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7527__A3 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__B2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4621__I _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8488__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A2 _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7153__B _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _0628_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5474__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8760_ _0159_ clknet_3_6_0_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ _1230_ _1473_ _1476_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7711_ _3002_ _2958_ _3075_ _2227_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_80_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4923_ _0470_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8691_ _0090_ clknet_leaf_42_wb_clk_i as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7642_ _3009_ _2993_ _2954_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4854_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4785_ _0317_ _0324_ _0345_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7573_ _1170_ _2849_ _2942_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8003__I _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6524_ _1973_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7151__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _0301_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7842__I _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6886__C _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5406_ _4186_ _0905_ _0907_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6386_ _1822_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8125_ _3425_ _3439_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5337_ _3935_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5362__I _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7454__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ as2650.r123\[0\]\[7\] as2650.r123_2\[0\]\[7\] _3886_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8056_ as2650.stack\[7\]\[5\] _3371_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7007_ _2366_ _2388_ _2403_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _0471_ _0637_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8403__A1 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7206__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7289__I _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6193__I _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6965__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _1684_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__A1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__I _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5940__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5153__B1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__B _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8069__B _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5456__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7701__B _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8583__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__B2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7420__C _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__I _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__A2 _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7381__A1 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6184__A2 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8731__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7381__B2 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4570_ _4064_ _4001_ _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6987__B _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7133__A1 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ _1310_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6171_ as2650.psl\[1\] _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5182__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5447__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5053_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5998__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8812_ _0211_ clknet_leaf_64_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4526__I _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8743_ _0142_ clknet_leaf_61_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5955_ _1464_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7837__I _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _4188_ _0428_ _0465_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_80_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8674_ _0073_ clknet_leaf_25_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5886_ _4006_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7625_ _2862_ _2989_ _2991_ _2610_ _2992_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4837_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6175__A2 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7556_ _0727_ _0669_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ _0285_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6507_ _0393_ _1951_ _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7124__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _3988_ _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7487_ _1151_ net9 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7675__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6438_ _1872_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5686__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6369_ _4011_ _1816_ _1817_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8108_ _1295_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8039_ _1494_ _2121_ _3365_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5820__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8604__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__C _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4661__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6938__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8754__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6953__A4 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5374__B1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A2 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7482__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7115__A1 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7666__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5677__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A1 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6826__I _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8091__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6929__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A1 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _4170_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5671_ _1187_ _1208_ _1209_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7410_ _0426_ _2633_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4622_ _4170_ _3959_ _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8390_ _3485_ _3694_ _3695_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7341_ _2668_ _2713_ _2714_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4553_ _4047_ _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7106__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__I _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4484_ _3953_ _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7272_ as2650.psu\[2\] _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5668__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ as2650.stack\[1\]\[2\] _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8627__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _4175_ _1102_ _1404_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4891__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5105_ as2650.r0\[6\] _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6085_ _1408_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6093__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _0456_ _0556_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__A2 _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__A1 _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6987_ _1573_ _2382_ _2383_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7593__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8726_ _0125_ clknet_leaf_27_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5938_ _1451_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4946__A3 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8657_ _0056_ clknet_leaf_32_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5869_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7608_ _1262_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7896__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8588_ _1739_ _2433_ _2576_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7539_ _2905_ _2908_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7648__A2 _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput12 net12 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 net23 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7820__A2 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4398__A1 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8533__B1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7639__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8257__B _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8064__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5460__I _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7811__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5822__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4625__A2 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6910_ _0359_ _0433_ _0564_ _2307_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_130_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7890_ _1380_ _1378_ _0911_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6841_ _1673_ _2246_ _2249_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7575__A1 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6505__B _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6291__I _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4389__A1 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _1913_ _2191_ _2195_ as2650.r123_2\[1\]\[1\] _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8511_ _1265_ _3797_ _3799_ _3800_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_50_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7327__B2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__S _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8442_ _3738_ _1946_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7878__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5654_ as2650.stack\[6\]\[8\] _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4605_ net10 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8373_ _3042_ _3406_ _3678_ _3412_ _1688_ _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5635__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6550__A2 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _0965_ _1127_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7324_ _2698_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4536_ _4043_ _4062_ _4115_ _4116_ _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _2630_ _2293_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ as2650.r0\[0\] _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5571__S _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6206_ _1142_ _1694_ _1697_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7186_ _2268_ _2564_ _1305_ _2424_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4398_ _3906_ _3978_ _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8055__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ _1632_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5370__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6068_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6369__A2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7566__A1 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__B2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8709_ _0108_ clknet_leaf_66_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7318__A1 _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7869__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7246__B _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5545__I _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8294__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6376__I _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7000__I _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4543__A1 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5370_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4321_ as2650.halted _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8285__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5099__A2 _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7493__B1 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ _0992_ _2398_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6835__A3 _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4846__A2 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8037__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8588__A3 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6599__A2 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _3260_ _1518_ _3294_ _3295_ _3296_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7873_ _3230_ _3210_ _3231_ _0903_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6824_ _1280_ net10 _1284_ _1289_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8815__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6755_ _1157_ _0982_ _1043_ _2171_ _2161_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7845__I _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _3971_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4782__B2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6686_ _2118_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8425_ _2353_ _3724_ _3727_ _2496_ _3728_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7315__A4 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7720__A1 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4534__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8356_ _3398_ _3660_ _3662_ _2569_ _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5568_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7307_ _2681_ _2227_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8276__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4519_ _4099_ _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8287_ _3589_ _3592_ _3596_ _2279_ _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_65_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5499_ _1007_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7513__C _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7238_ _2613_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7169_ _2358_ _2546_ _2550_ _2280_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7787__A1 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__I as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7711__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8586__I _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8267__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A1 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__I _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8019__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__A1 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8838__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _0430_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5005__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7950__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5556__A3 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7950__B2 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ _4260_ _1845_ _1992_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4764__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6502__C _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6471_ _1923_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6505__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7702__B2 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _3520_ _3521_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5422_ _0916_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5118__C _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8141_ _3390_ _3454_ _3455_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8258__A2 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5353_ _4120_ _0897_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6269__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4304_ _3884_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6269__B2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8072_ _3387_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7333__C _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5284_ _0812_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_82_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7023_ _1645_ _1503_ _1625_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__S _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__A1 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _1318_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7856_ _3160_ _4251_ _1567_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8194__A1 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _3917_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7787_ _2661_ _3137_ _3146_ _3148_ _3011_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4999_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6738_ _1912_ _2164_ _2169_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5095__I _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8497__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6669_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8408_ net39 _3654_ _3655_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7524__B _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8339_ _2470_ _3505_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6654__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8421__A2 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A2 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4994__B2 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8185__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7932__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8488__A2 _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__I _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A3 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__C _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7448__B1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7463__A3 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8660__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ as2650.stack\[1\]\[13\] _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6974__A2 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7710_ as2650.addr_buff\[0\] as2650.addr_buff\[1\] as2650.addr_buff\[2\] _3075_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4922_ _0483_ _0328_ _0346_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4985__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8690_ _0089_ clknet_leaf_39_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8176__A1 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7641_ _2617_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4853_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7923__A1 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _2896_ _2941_ _2847_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4784_ _4292_ _0346_ _4284_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6523_ _1975_ _1976_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _1832_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7151__A2 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5405_ _4185_ _0893_ _0961_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5162__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _1841_ _1548_ _4161_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5162__B2 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8124_ _4272_ _3427_ _3430_ _3432_ _3438_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_115_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _0892_ _4034_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8100__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8055_ _2130_ _3369_ _3374_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5267_ as2650.r0\[2\] _0572_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7006_ _2388_ _2401_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6662__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _0754_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6965__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7908_ _0564_ _1721_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4976__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8167__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8167__B2 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7839_ _3172_ _3197_ _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6717__A2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5153__A1 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8069__C _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8683__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7701__C _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__I _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5208__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__B2 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8158__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6169__B1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7905__A1 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6708__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6184__A3 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5144__A1 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ _4108_ _4069_ _0424_ _1661_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ _0382_ _0639_ _0649_ _4059_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5052_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4655__B1 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4807__I _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8811_ _0210_ clknet_leaf_64_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8742_ _0141_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5954_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4905_ _0462_ _4188_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8673_ _0072_ clknet_leaf_25_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5885_ _1391_ _1406_ _1407_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_139_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7624_ _1255_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4836_ as2650.r123\[0\]\[2\] as2650.r123_2\[0\]\[2\] as2650.psl\[4\] _0399_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7555_ _0656_ _0577_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4767_ _0325_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6506_ _0386_ _1815_ _1857_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7486_ as2650.pc\[4\] _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7124__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8321__A1 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _4237_ _4244_ _4249_ _4276_ _4277_ _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6437_ _1876_ _1879_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_122_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6883__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6368_ _1821_ _1823_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8107_ _3421_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ _3943_ _3990_ _0866_ _0863_ _4018_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6299_ as2650.stack\[3\]\[10\] _1759_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6635__A1 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7832__B1 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8038_ as2650.stack\[4\]\[12\] _3361_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5322__B _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8388__A1 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6938__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7060__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8560__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8312__A1 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7115__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6874__A1 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7003__I _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8379__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__A3 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6929__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6842__I _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6063__B _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__I _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_32_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5670_ as2650.stack\[6\]\[10\] _1202_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8551__A1 _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _4201_ _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _1128_ _4268_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4552_ _4117_ _4132_ _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8303__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7106__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7271_ _2644_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ _4063_ _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6222_ _1463_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5668__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4340__A2 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6153_ _1397_ _1405_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6617__A1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5104_ _0658_ _0562_ _4073_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6084_ _1546_ _1579_ _1275_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__A2 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5035_ _4114_ _0589_ _0595_ _4277_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__A3 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7042__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6986_ _1087_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5937_ _1193_ _1450_ _1453_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8725_ _0124_ clknet_leaf_24_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5368__I _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8656_ _0055_ clknet_leaf_31_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5868_ _3934_ _1245_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7345__A2 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8542__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7607_ _0976_ _2971_ _2973_ _2975_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4819_ _4060_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8587_ _1739_ _2441_ _3870_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5799_ _1325_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7538_ _2855_ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7516__C _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5108__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7469_ as2650.stack\[2\]\[4\] _0939_ _2797_ as2650.stack\[3\]\[4\] _2840_ _2841_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_107_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput13 net49 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput24 net24 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7281__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__B2 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A2 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7584__A2 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8871__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4398__A2 _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7336__A2 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8533__B2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5898__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__A2 _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6847__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6311__A3 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__I _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__B _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4357__I _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__A3 _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__A1 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8221__B1 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6840_ _2247_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2192_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4389__A2 _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8510_ _1591_ _1417_ _3175_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5722_ _1243_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8524__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7327__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8441_ _0303_ _3733_ _3740_ _3742_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5338__A1 _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8499__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _1186_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4820__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _4039_ _4133_ _4184_ _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8372_ _3132_ _3050_ _3408_ _3677_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5584_ _1130_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ _0950_ as2650.stack\[7\]\[1\] as2650.stack\[6\]\[1\] _0939_ _0972_ _2698_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4535_ _3980_ _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7254_ as2650.addr_buff\[0\] _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4466_ _4044_ _4046_ _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6205_ as2650.stack\[0\]\[2\] _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8744__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5510__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ _2486_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4397_ _3976_ _3977_ _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8167__C _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4695__C _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6136_ _3903_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A2 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _1372_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5018_ as2650.r0\[5\] _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5098__I _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6969_ net25 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8708_ _0107_ clknet_leaf_22_wb_clk_i as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8515__A1 _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5329__A1 _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8639_ _0038_ clknet_leaf_3_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6829__A1 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4886__B _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5804__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5002__S _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A2 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8506__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8617__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4543__A2 _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5740__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _3900_ _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7493__B2 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7941_ _1524_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__I _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7872_ _2648_ _1387_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _1278_ _2226_ _2230_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5559__A1 _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6220__A2 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ as2650.r123_2\[0\]\[5\] _2154_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _3995_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6685_ _1154_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4550__I _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8424_ _1221_ _3421_ _3388_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5636_ _1176_ _1177_ _1076_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7720__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8355_ _2252_ _3661_ _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5567_ as2650.pc\[0\] _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5731__A1 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7861__I _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7306_ as2650.addr_buff\[1\] _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4518_ _4080_ _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8286_ _1168_ _3405_ _3595_ _2720_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5498_ _1009_ as2650.stack\[5\]\[14\] as2650.stack\[4\]\[14\] _0946_ _1049_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_137_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7484__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _0437_ _1713_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6287__A2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ _3963_ _4029_ _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7168_ _2377_ _2531_ _2542_ _2548_ _2549_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7236__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _1257_ _0898_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7099_ _2483_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7787__A2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5798__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7101__I _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4470__A1 as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8360__C _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7711__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7227__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4836__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7778__A2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__I0 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4635__I _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8107__I _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7011__I _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6202__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7950__A2 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4764__A2 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _0821_ _1881_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8140_ net52 _3418_ _3321_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5352_ _4187_ _0905_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4303_ _3883_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7466__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6269__A2 _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8071_ _2311_ _3386_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7466__B2 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5283_ _0815_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ _3976_ _2412_ _2416_ _2415_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__B _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4545__I _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7924_ _3153_ _0654_ _2481_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__A1 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6729__B1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7855_ _2156_ _2704_ _3214_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8194__A2 _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6806_ _2215_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4998_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7786_ _2661_ _3147_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6737_ as2650.r123_2\[0\]\[1\] _2165_ _2168_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5952__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6668_ _1079_ _1184_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8407_ _3696_ _3486_ _3707_ _3453_ _3711_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5619_ _1157_ _1158_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5704__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6599_ _0667_ _2050_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8338_ _2300_ _1525_ _3641_ _3645_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_2_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5180__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8269_ _3574_ _3578_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6000__I _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7209__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6680__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7224__A4 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6432__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__I _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A3 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8371__B _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__A2 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6670__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7393__B1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7932__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7696__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7448__A1 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7448__B2 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7999__A2 _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8805__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6066__B _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__I _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__A1 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _1466_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4921_ _0320_ _0338_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7676__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8176__A2 _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7640_ _0956_ _2800_ _2993_ _3006_ _3007_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4852_ as2650.r0\[4\] _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7923__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7571_ _2901_ _2912_ _2940_ _2845_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4783_ _0321_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _0666_ _0573_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8479__A3 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _4236_ _1837_ _1907_ _1908_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ as2650.r123\[0\]\[0\] _0909_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _4095_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5162__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7439__A1 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8123_ _3433_ _3435_ _3437_ _3397_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5335_ _0569_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8100__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8054_ as2650.stack\[7\]\[4\] _3371_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6111__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5266_ as2650.r0\[1\] _0785_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4984__B _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7005_ _1632_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _0755_ _0635_ _0628_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A1 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6414__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__B2 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6965__A3 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7907_ _3260_ _0548_ _1525_ _3263_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8167__A2 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4440__A4 _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ _1849_ _3198_ _1622_ _0872_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7914__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4728__A2 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7769_ _2629_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5834__I _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5153__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8828__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7602__A1 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6169__B2 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7905__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7669__A1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7669__B2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5744__I _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5120_ _0381_ _0651_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8094__A1 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5051_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4655__A1 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4655__B2 _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8810_ _0209_ clknet_leaf_64_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4407__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8741_ _0140_ clknet_leaf_62_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _1112_ _1447_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _3937_ _0428_ _0463_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5884_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8672_ _0071_ clknet_leaf_24_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _1188_ _2990_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4835_ _4245_ _0307_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5907__A1 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7554_ _2917_ _2923_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _0324_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6580__A1 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6505_ _0374_ _1808_ _1815_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7485_ _2854_ _2855_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _4125_ _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6332__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6436_ _1883_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6332__B2 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6883__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _3975_ _3979_ _1813_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_103_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8106_ _3420_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5318_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6298_ _1487_ _1755_ _1760_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7832__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _4035_ _0771_ _0807_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8037_ _1492_ _3359_ _3364_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7832__B2 _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8388__A2 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__A1 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7060__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8560__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8650__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4889__B _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7265__B _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__A1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5429__A3 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8379__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4652__A4 _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8000__A1 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _4200_ _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6562__A1 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4551_ _4126_ _4131_ _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8303__A2 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7270_ _2645_ as2650.stack\[5\]\[0\] as2650.stack\[4\]\[0\] _1008_ _2646_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4482_ _4050_ _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5117__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _1134_ _1704_ _1705_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8067__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _0874_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _4071_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7814__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _1103_ _0436_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4628__A1 _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _4042_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7042__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6985_ _1286_ _2235_ _3985_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5649__I _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8724_ _0123_ clknet_leaf_46_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5936_ as2650.stack\[0\]\[8\] _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8673__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8655_ _0054_ clknet_leaf_22_wb_clk_i as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5867_ _1385_ _1388_ _1390_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__8542__A2 _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7606_ _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4818_ _4058_ _3919_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8586_ _3869_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ _0872_ _1329_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7537_ _2906_ _2854_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4749_ _0309_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5384__I _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6305__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__A2 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7468_ _2644_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net14 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput25 net25 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _0665_ _0505_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput36 net36 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7399_ _2723_ _2758_ _2765_ _2724_ _2771_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6608__A2 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7805__A1 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A4 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7033__A2 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5044__A1 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__B _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7336__A3 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8533__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5898__A3 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4638__I _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6853__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8696__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8221__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8221__B2 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A1 _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4373__I _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6783__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6770_ _2189_ _2194_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5721_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8440_ as2650.r123\[2\]\[1\] _3741_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5338__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _4039_ _4183_ _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8371_ _2876_ _3676_ _3060_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5583_ _1125_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8288__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4534_ _4064_ _4066_ _4113_ _4114_ _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7322_ _2695_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8288__B2 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7253_ _2337_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4465_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _4045_ _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6204_ _1448_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7184_ _2442_ _3916_ _2515_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7352__C _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4396_ as2650.idx_ctrl\[0\] _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5510__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _1526_ _1572_ _1621_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6066_ _1557_ _1560_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__I _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5017_ _4099_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7015__A2 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8212__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8212__B2 _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6968_ net49 _2352_ _2365_ _1438_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8707_ _0106_ clknet_leaf_24_wb_clk_i as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5919_ _1441_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6899_ _1570_ _1259_ _1602_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8638_ _0037_ clknet_leaf_3_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6526__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8569_ _3850_ _3855_ _4036_ _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8279__A1 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__I _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6829__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4458__I _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8451__A1 _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__I _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8203__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5017__A1 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6765__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8506__A2 _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7190__A1 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4543__A3 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5740__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6848__I _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__I _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7493__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6069__B _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8442__A1 _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6583__I _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _3205_ _0722_ _2547_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7871_ as2650.overflow _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6822_ _1104_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5559__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _2072_ _2151_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ _1194_ _1237_ _1238_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7347__C _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6684_ _2128_ _2119_ _2129_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8423_ _1221_ _3647_ _3726_ _2371_ _3106_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5635_ as2650.pc\[7\] _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8354_ _3001_ _3626_ _3628_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5731__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7305_ _4271_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4517_ _4097_ _3896_ _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8285_ _2777_ _2910_ _3506_ _3594_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5497_ _0741_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7484__A2 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7236_ _1117_ _4069_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _4025_ _3900_ _4028_ _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7167_ _1741_ _2283_ _2389_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4379_ _3957_ _3959_ _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7236__A2 _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6118_ _1260_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7810__C _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7098_ _1302_ _2404_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8194__B _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ _1534_ _1542_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5798__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6747__A1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4741__I _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4525__A3 _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5572__I _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__C _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__B2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8424__A1 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5238__B2 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5789__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4836__I1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6738__A1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5747__I _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8734__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__I _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5961__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7163__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8884__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6910__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4302_ _3882_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8070_ _2339_ _2589_ _3382_ _3385_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5282_ _0818_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _2265_ _2400_ _2412_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7911__B _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6977__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7923_ _3205_ _0682_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__A2 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7854_ _0308_ _3162_ _3212_ _3213_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6729__B2 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7926__B1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ as2650.r123\[3\]\[7\] _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5657__I _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7785_ _1054_ _2654_ _3137_ _2271_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4997_ net9 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5401__A1 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6736_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5952__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7154__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _1120_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7154__B2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8406_ _2863_ _3083_ _3709_ _2389_ _3710_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5618_ _1160_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5704__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _1792_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8337_ _2983_ _3642_ _3644_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5549_ as2650.cycle\[3\] _1088_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5392__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8268_ _3576_ _3549_ _3577_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_117_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5468__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7219_ _4122_ _2594_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8199_ _2757_ _3486_ _3511_ _3452_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8607__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8406__A1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7209__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8406__B2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7112__I _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8757__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4672__S _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A4 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7393__A1 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5567__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7448__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5459__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__B2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8118__I _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6959__A1 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7957__I as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ _4291_ _4156_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _4099_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7570_ _2623_ _2913_ _2911_ _2932_ _2939_ _2654_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_4782_ _0330_ _0342_ _0343_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _1972_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7136__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7625__C _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _4244_ _1835_ _1837_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5403_ _0909_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6383_ _4214_ _1839_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8122_ _4272_ _3436_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4370__A1 _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5334_ _0496_ _0843_ _0891_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8053_ _2128_ _3369_ _3373_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5265_ _0820_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _1718_ _2399_ _2400_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ _0627_ _0585_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4673__A2 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A3 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8472__B _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7867__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7906_ _3260_ _3261_ _3262_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7837_ _2231_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7375__A1 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7768_ _1254_ _0437_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _1860_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7127__A1 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7699_ _3053_ _3055_ _3064_ _1735_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_109_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5689__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__A2 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6946__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5850__I _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5310__C2 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A3 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7366__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4719__A3 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__A2 _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5050_ as2650.r123\[0\]\[4\] as2650.r123_2\[0\]\[4\] as2650.psl\[4\] _0611_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5852__A1 _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__I as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7687__I _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4407__A2 _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8740_ _0139_ clknet_leaf_44_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5952_ _1237_ _1458_ _1462_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4903_ _0363_ _0368_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8671_ _0070_ clknet_leaf_78_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7357__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5883_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7622_ _1177_ _2897_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4834_ _0373_ _4220_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5000__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7553_ _2816_ _2910_ _2922_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _0326_ _0289_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5935__I _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _0350_ _1952_ _1957_ _1958_ _1807_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7484_ _1159_ _1652_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _4250_ _4251_ _4275_ _4067_ _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_101_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6435_ _1886_ _1890_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8105_ _1622_ _2287_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7371__B _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6766__I _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8085__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6297_ as2650.stack\[3\]\[9\] _1759_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6096__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8036_ as2650.stack\[4\]\[11\] _3361_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7832__A2 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ as2650.r123\[1\]\[6\] _0600_ _0806_ _0408_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_76_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5179_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7596__A1 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7348__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8869_ _0268_ clknet_leaf_66_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6006__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4582__A1 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7520__B2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4334__A1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8808__D _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__A2 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7823__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__A1 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6929__A4 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8000__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4550_ _4130_ _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _4061_ _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ as2650.stack\[1\]\[1\] _1475_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4325__A1 _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8067__A2 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6151_ _0869_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _0585_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ _0538_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7814__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__A1 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5033_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7578__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6984_ _1609_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8818__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6250__A1 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8723_ _0122_ clknet_leaf_46_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4800__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8654_ _0053_ clknet_leaf_24_wb_clk_i as2650.stack\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5866_ _4009_ _0851_ _1391_ _0899_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6002__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7605_ _2648_ as2650.stack\[7\]\[7\] as2650.stack\[6\]\[7\] _1006_ _0953_ _2974_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0378_ _4231_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8585_ _4191_ _1383_ _3851_ _3868_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__5665__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6553__A2 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _4064_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7536_ as2650.pc\[4\] _0558_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4564__A1 _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4748_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7467_ _2645_ as2650.stack\[1\]\[4\] as2650.stack\[0\]\[4\] _1008_ _2839_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6305__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _4253_ _4258_ _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4316__A1 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6418_ _1788_ _1873_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput15 net15 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput26 net26 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ _2259_ _2228_ _2770_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput37 net37 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6496__I _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8058__A2 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _3936_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__A1 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5816__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8019_ _3350_ _1208_ _3354_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6445__B _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7569__B2 _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7120__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5044__A2 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8297__A2 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5504__B1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5016__S _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__I _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8126__I _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8221__A2 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6232__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6783__A2 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5720_ _1103_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4794__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7186__B _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5651_ _1190_ _1076_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5485__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7732__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ _4182_ _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8370_ net38 _3675_ _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5418__C _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5582_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7321_ _1037_ as2650.stack\[5\]\[1\] as2650.stack\[4\]\[1\] _1009_ _2696_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _4041_ _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7914__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8288__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _2360_ _1395_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4464_ _3887_ _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6203_ _1134_ _1694_ _1695_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7183_ _2558_ _2561_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4395_ as2650.idx_ctrl\[1\] _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _1623_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _4020_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5016_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _0411_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8640__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _2353_ _2364_ _2352_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8480__B _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8790__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5918_ as2650.r123_2\[3\]\[2\] _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4785__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8706_ _0105_ clknet_leaf_34_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ _2281_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8637_ _0036_ clknet_leaf_3_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5849_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6526__A2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _3854_ _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7519_ _0949_ as2650.stack\[7\]\[5\] as2650.stack\[6\]\[5\] _0921_ _0952_ _2890_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8279__A2 _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8499_ _0439_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8451__A2 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4474__I _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8203__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5017__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6765__A2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7962__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7962__B2 _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7714__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__I _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__C _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8663__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8442__A2 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6453__A1 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4384__I _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7870_ _3207_ _0349_ _3226_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6821_ _2228_ _2229_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7953__A1 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ _2041_ _2164_ _2180_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ as2650.stack\[6\]\[14\] _1231_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6683_ as2650.stack\[4\]\[3\] _2124_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8422_ _2261_ _2481_ _3725_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5634_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8353_ _2252_ _3659_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5192__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5565_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5731__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7304_ _1089_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7469__B1 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4516_ _4096_ _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8284_ _2920_ _3593_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5496_ as2650.r123\[0\]\[6\] _0962_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_137_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7235_ _2610_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4559__I _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4447_ _4026_ _4027_ _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6692__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7166_ _2547_ _1099_ _2377_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4378_ _3958_ _3944_ _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6117_ _1611_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6774__I _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _2457_ _4118_ _2481_ _2376_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8197__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7999_ as2650.stack\[6\]\[2\] _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7944__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6904__C1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5183__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7273__C _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8686__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7227__A3 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8424__A2 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7632__B1 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A3 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7935__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7448__C _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7163__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8360__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5174__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5763__I _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6910__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8279__C _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _0906_ _4209_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4921__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4301_ as2650.ins_reg\[0\] _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_126_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5281_ _0830_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _3977_ _2412_ _2413_ _2415_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5477__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6674__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8415__A2 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6426__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__A2 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7922_ _3264_ _3277_ _3278_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7853_ _1563_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6729__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7926__A1 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5938__I _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6804_ _2214_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7784_ _3138_ _3145_ _2528_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4996_ _0417_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5401__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _2157_ _0981_ _2160_ _0310_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _2061_ _2103_ _2115_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8405_ _3696_ _3567_ _2664_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5617_ _1125_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5165__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6597_ _2015_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8336_ _3588_ _3643_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4912__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5548_ as2650.cycle\[2\] _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8103__A1 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_opt_3_0_wb_clk_i clknet_3_1_0_wb_clk_i clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8267_ _3575_ _0681_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5479_ _1025_ _0966_ _1031_ _0982_ _0983_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_132_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7218_ _2221_ _2531_ _1106_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7862__B1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8198_ _1145_ _3274_ _3226_ _3504_ _3510_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7149_ _2530_ _2519_ _2531_ _2362_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8406__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6417__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6968__A2 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7090__A1 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__S0 _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4979__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7393__A2 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8590__B2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout50 net37 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8342__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8342__B2 _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6679__I _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4927__I _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7303__I _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__B1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8701__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8562__C _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5631__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7908__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8581__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8851__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A1 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ _4172_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _0579_ _0786_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8333__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7136__A2 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _4246_ _1853_ _1900_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6895__A1 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _4215_ _0914_ _0956_ _0957_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6382_ _1838_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8121_ _4123_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5333_ as2650.r123\[1\]\[7\] _0600_ _0890_ _4210_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4370__A2 _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6647__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ as2650.stack\[7\]\[3\] _3371_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5264_ _0796_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _2299_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4837__I _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5195_ _0750_ _0751_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8472__C _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7905_ _2570_ _0594_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7836_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7767_ _2506_ _3128_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4979_ _0538_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6718_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7127__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7698_ _3059_ _3063_ _2467_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _2080_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5109__S _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6886__A1 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__A3 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8319_ _0875_ _0885_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6638__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8724__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5310__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5310__B2 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6962__I _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8874__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4482__I _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8563__A1 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4352__A2 _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4657__I _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5301__A1 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5852__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5604__A2 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ as2650.stack\[0\]\[14\] _1460_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ as2650.holding_reg\[3\] _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8670_ _0069_ clknet_3_2_0_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5882_ _3956_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8554__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7621_ _2983_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4833_ _0316_ _0349_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_61_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7552_ _2918_ _2913_ _2921_ _2635_ _2219_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _4285_ _4262_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8306__A1 _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _0370_ _1850_ _1823_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7483_ _2853_ net1 _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4695_ _4032_ _4261_ _4274_ _4111_ _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6868__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6434_ _1887_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5540__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8747__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__A2 _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _4014_ _3964_ _4019_ _1818_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8104_ _3390_ _3417_ _3419_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ net3 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _1756_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7293__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _1490_ _3359_ _3363_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6096__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _0774_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5178_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8868_ _0267_ clknet_leaf_65_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7348__A2 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8545__A1 _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7819_ _3994_ _1065_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8799_ _0198_ clknet_leaf_19_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__I _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6022__I _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7562__B _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6957__I _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5531__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__I _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__A2 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7339__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8536__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6641__B _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8412__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7028__I _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4480_ _4055_ _4060_ _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4325__A2 _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6150_ _1599_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _4264_ _0552_ _0650_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__7275__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6078__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4387__I _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1576_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7814__A3 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _4239_ _0550_ _0590_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6816__B _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__B1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7578__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5589__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _2375_ _2376_ _2377_ _2379_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6250__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8722_ _0121_ clknet_leaf_46_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _1448_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5865_ _1083_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8653_ _0052_ clknet_leaf_35_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _2695_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4816_ _0378_ _4229_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _1328_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8584_ _3885_ _2329_ _3761_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7535_ _2859_ _2856_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4747_ _0310_ _4223_ _0308_ _4215_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7466_ _0950_ as2650.stack\[7\]\[4\] as2650.stack\[6\]\[4\] _0939_ _0972_ _2838_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_135_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4678_ _4256_ _3894_ _4087_ _4257_ _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6417_ _1787_ _1790_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4316__A2 _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _2217_ _2769_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput16 net16 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput38 net38 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ _1771_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7266__A1 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6279_ as2650.stack\[2\]\[3\] _1746_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8018_ as2650.stack\[5\]\[10\] _3352_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8518__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8388__B _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5504__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4935__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8221__A3 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8509__A1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7980__A2 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__A2 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5766__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8142__I _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7186__C _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _4223_ _1126_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _4142_ _4147_ _4153_ _4181_ _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5743__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7320_ _2643_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4532_ _4067_ _4112_ _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7496__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7251_ _1673_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6299__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4463_ _3891_ as2650.ins_reg\[1\] _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ as2650.stack\[0\]\[1\] _1460_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7182_ _2539_ _2560_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4394_ _3971_ _3974_ _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7248__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _1627_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _4202_ _1430_ _1406_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__I _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5015_ _0568_ _0571_ _0574_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7420__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7420__B2 _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ _2355_ _2359_ _2363_ _1577_ _2275_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_74_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8705_ _0104_ clknet_leaf_32_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5917_ _1440_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6897_ _1262_ _2292_ _2294_ _2295_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_107_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8636_ _0035_ clknet_leaf_2_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _1273_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8567_ _1393_ _1589_ _3853_ _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5779_ _1292_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_120_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7518_ _2643_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8498_ _0968_ _3786_ _3788_ _3624_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7487__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7449_ _2816_ _2811_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7239__A1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7131__I _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__C _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7411__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5586__I _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__I _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5725__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__A2 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8808__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8137__I _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__I _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7041__I _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6880__I _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6205__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ _1713_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7197__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ as2650.r123_2\[0\]\[4\] _2165_ _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5964__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5702_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6682_ _1147_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8421_ _3563_ _3718_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5633_ _0870_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8352_ _3001_ _3631_ _3632_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7644__C _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ _1079_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7303_ _1409_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4515_ as2650.r0\[7\] _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7469__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8283_ _2228_ _3573_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _1046_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7234_ _2219_ _1733_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4446_ _3996_ _3949_ _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7165_ _1269_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6692__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4377_ _3899_ _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6116_ _3972_ _1088_ _3973_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7096_ _2462_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5180__B _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4575__I _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6047_ _0876_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8491__B _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _1185_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6949_ _2341_ _2343_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8619_ _0018_ clknet_leaf_25_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6904__B1 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6904__C2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5183__A2 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6132__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7880__A1 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7062__S _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4694__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4485__I _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7632__A1 _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A2 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7632__B2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5789__A4 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7796__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7935__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4749__A2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A1 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7163__A3 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8360__A2 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6371__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8630__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6910__A3 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__A2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4300_ net26 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5280_ _0832_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6123__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8780__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6426__A2 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4437__A1 _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7921_ _1350_ _3240_ _3040_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _1666_ _1388_ _3211_ _1389_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7926__A2 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6803_ as2650.r123\[3\]\[6\] _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5937__A1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7783_ _3141_ _3144_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6734_ _2153_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6665_ as2650.r123_2\[2\]\[7\] _1948_ _2114_ _2043_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8404_ _3696_ _2297_ _3562_ _3708_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5616_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6596_ _2047_ _2020_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8335_ _2983_ _3642_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5547_ _3912_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4912__A2 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8103__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6114__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5478_ _1027_ _1028_ _1030_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8266_ _3575_ _0681_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_133_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7217_ _2158_ _1609_ _2590_ _2592_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__6665__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7862__A1 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _4006_ _4009_ _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__7862__B2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8197_ _1720_ _3509_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7148_ _1093_ _1089_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7079_ _2268_ _2460_ _2372_ _2463_ _2383_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7090__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__S1 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4979__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout51 net33 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8653__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8342__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6353__A1 _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4903__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6105__A1 _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7302__B1 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6408__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7605__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__B2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4943__I _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7908__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8030__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4780_ _4154_ _0322_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_35_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8333__A2 _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5147__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _1853_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7541__B1 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5401_ _4197_ _0904_ _0894_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6895__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _4003_ _1503_ _3951_ _1810_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_103_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8097__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8120_ _2251_ _4236_ _3434_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5332_ _0316_ _0862_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_126_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6647__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5263_ as2650.r0\[5\] _0399_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8051_ _2126_ _3369_ _3372_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4658__A1 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6538__C _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7002_ _1741_ _2389_ _2396_ _2398_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5194_ as2650.holding_reg\[6\] _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5083__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4853__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7904_ _3153_ _0556_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8884_ _0283_ clknet_leaf_41_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8676__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8021__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7835_ _3173_ _3183_ _3187_ _3195_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_93_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7766_ _1043_ _2977_ _3123_ _2665_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4978_ _0521_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6717_ _0906_ _1827_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_138_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _2816_ _3050_ _3051_ _2379_ _3062_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_137_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8324__A2 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6648_ _2077_ _2081_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5138__A2 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _0564_ _1846_ _1956_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8088__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4897__B2 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8318_ _3574_ _3578_ _3625_ _3602_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7832__C _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8249_ _3441_ _3559_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7404__I _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5310__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8260__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__I _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4821__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__A2 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6326__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6877__A2 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4888__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8079__A1 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7826__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8699__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7189__C _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5950_ _1230_ _1458_ _1461_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4812__A1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _0462_ _3937_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7984__I _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5881_ _1253_ _1375_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8554__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7620_ _2909_ _2985_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_61_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4832_ _4281_ _0388_ _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7762__B1 _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7551_ _2919_ _2920_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4763_ _4285_ _4262_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _1953_ _1846_ _1955_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7482_ as2650.pc\[5\] _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4694_ _4072_ _4267_ _4273_ _4079_ _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6868__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _1884_ _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6364_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5540__A2 _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8103_ _3400_ _3418_ _3321_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7817__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4848__I _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ _4095_ _0872_ _4109_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_130_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6295_ _1478_ _1755_ _1758_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7293__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8490__A1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8034_ as2650.stack\[4\]\[10\] _3361_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5246_ _0777_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5177_ _4098_ _4102_ _4105_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8242__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4583__I _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8867_ _0266_ clknet_leaf_65_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8545__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7818_ _1527_ _2288_ _1580_ _3178_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8798_ _0197_ clknet_leaf_19_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7749_ _2676_ _3105_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6303__I _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6308__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7843__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7562__C _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5531__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5082__C _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8481__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8841__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5295__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7036__A2 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__I _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8536__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5770__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__B _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _3944_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _1575_ _1260_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8472__A1 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7814__A4 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _0591_ _0543_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4628__A4 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__B2 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _2378_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5589__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8721_ _0120_ clknet_leaf_29_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5933_ _1449_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_50_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8527__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8652_ _0051_ clknet_leaf_32_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5864_ _4196_ _1389_ _1074_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7603_ _1037_ as2650.stack\[5\]\[7\] as2650.stack\[4\]\[7\] _0942_ _2972_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4815_ _4259_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8583_ net27 _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8714__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5210__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7534_ _2903_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4746_ _4246_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5761__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7465_ _2695_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4677_ as2650.r123\[1\]\[2\] as2650.r123\[0\]\[2\] as2650.r123_2\[1\]\[2\] as2650.r123_2\[0\]\[2\]
+ _3891_ _4045_ _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6416_ _1784_ _1800_ _1871_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8864__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7396_ _0427_ _2390_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput17 net17 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput28 net28 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6347_ _1773_ _1775_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7266__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6278_ _1142_ _1744_ _1747_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5277__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7889__I _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8017_ _3350_ _1201_ _3353_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5229_ _0572_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6777__A1 _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5044__A4 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8518__A2 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6033__I _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__C1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4488__I _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7009__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7965__B1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8737__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8509__A2 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7193__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _4157_ _4158_ _4180_ _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5743__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6940__A1 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ as2650.pc\[1\] _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6878__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _4078_ _4094_ _4110_ _4111_ _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7496__A2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7250_ _2461_ _4046_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4462_ _4042_ _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6201_ _1451_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4393_ _3972_ _3911_ _3973_ _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7181_ as2650.cycle\[5\] _2553_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7248__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8445__A1 _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _1553_ _1615_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _0892_ _1540_ _1558_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _3884_ _3892_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6759__A1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__B _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _2362_ _1264_ _2358_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5957__I _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4861__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8704_ _0103_ clknet_leaf_33_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5916_ as2650.r123_2\[3\]\[1\] _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _3972_ _1286_ _1577_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8635_ _0034_ clknet_leaf_2_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7184__A1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _1372_ _4029_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8566_ _1378_ _1396_ _3851_ _3852_ _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5778_ _1311_ _1090_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6931__A1 _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__B _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7517_ _0944_ as2650.stack\[5\]\[5\] as2650.stack\[4\]\[5\] _0941_ _2888_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4729_ _4160_ _0290_ _0291_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8497_ _0968_ _3070_ _2426_ _3787_ _3786_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_68_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7448_ _2817_ _2521_ _2675_ _2807_ _2819_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7487__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5498__A1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5498__B2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ _2665_ _2712_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7239__A2 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8436__A1 _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4473__A2 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5670__A1 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7411__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4856__S0 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6922__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__I _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5551__B _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__I _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__B2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__I _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _2178_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5964__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _1233_ _1211_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7166__A1 _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _2126_ _2119_ _2127_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7992__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8420_ _2544_ _3715_ _3723_ _3155_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_31_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ _1150_ _1173_ _1174_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6913__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A2 _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8351_ _3018_ _3657_ _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5563_ _1080_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7302_ _2675_ _2662_ _2671_ _2676_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7469__A2 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ as2650.psl\[3\] _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8282_ _3443_ _3591_ _3281_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5494_ _1035_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7233_ _1117_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4445_ as2650.ins_reg\[5\] _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8418__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7164_ _2542_ _2543_ _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4376_ as2650.ins_reg\[2\] _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6115_ _1088_ _1294_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8328__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7095_ _2457_ _1736_ _2479_ _2292_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7232__I _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__B1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _1535_ _1427_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ _2123_ _3339_ _3341_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5687__I _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4591__I _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _2345_ _2231_ _2239_ _2292_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_81_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6879_ _2279_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8618_ _0017_ clknet_leaf_25_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6904__A1 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6904__B2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8549_ _3809_ _3837_ _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__A2 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8409__A1 _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7880__A2 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4694__A2 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7396__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4715__B _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6199__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5946__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7148__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6371__A2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6123__A2 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4685__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__I _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7052__I _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7623__A2 _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4437__A2 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7920_ _3265_ _3276_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7851_ _0978_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7387__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6802_ _2213_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7782_ _3053_ _2919_ _3143_ _2946_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4994_ _0549_ _0421_ _0550_ _4233_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5937__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6733_ _2154_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7936__B _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7139__A1 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6664_ _1770_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8403_ _3563_ _3704_ _3084_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5615_ as2650.pc\[5\] _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6595_ _2017_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8334_ _2984_ _3590_ _2986_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5546_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8265_ _0656_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5970__I _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _0977_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6114__A2 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7216_ _2591_ _2332_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4428_ _4008_ _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8196_ _2946_ _2765_ _3505_ _1145_ _3508_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7862__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7147_ _2372_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4359_ _3939_ _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _2456_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8575__B1 _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__I _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net29 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7565__C _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7550__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6353__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6041__I _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__A1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__I _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6105__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7302__B2 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__A1 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5092__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8030__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xwrapped_as2650_90 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7541__A1 _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _0913_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6380_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8587__B _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5331_ _4126_ _0868_ _0888_ _4282_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8050_ as2650.stack\[7\]\[2\] _3371_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5262_ as2650.r0\[6\] _0305_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5855__A1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7001_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4658__A2 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _0750_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6280__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout50_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7903_ _2471_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8883_ _0282_ clknet_leaf_40_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6126__I _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8021__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7834_ _1806_ _3188_ _3190_ _1313_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_63_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__B _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7765_ _2618_ _3123_ _3126_ _2362_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_71_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4977_ _4154_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7780__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ _2138_ _1757_ _2149_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7696_ _2217_ _3061_ _0438_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5186__B _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ _2074_ _2082_ _2097_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _0560_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8317_ _0875_ _0885_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8088__A2 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _1068_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6099__A1 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _3402_ _3546_ _3558_ _3425_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7835__A2 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8179_ _3466_ _3490_ _3491_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7599__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8260__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8620__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4821__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7771__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8251__I _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6326__A2 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7523__A1 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7523__B2 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4888__A2 _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7826__A2 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6655__B _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6262__A1 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ as2650.holding_reg\[3\] _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5880_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _4116_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7762__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__B _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7550_ _1539_ _2390_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4576__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _4160_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6501_ _4003_ _4030_ _1810_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_7481_ _2618_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4693_ _4272_ _3967_ _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7514__A1 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7514__B2 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ as2650.r0\[3\] _0785_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4879__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6363_ _3962_ _3965_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7505__I _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8102_ _3388_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5314_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7817__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6294_ as2650.stack\[3\]\[8\] _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5828__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8033_ _1487_ _3359_ _3362_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _0780_ _0803_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5025__I _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8490__A2 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8643__CLK clknet_opt_2_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ _0730_ _4072_ _4074_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4864__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8242__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8793__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8866_ _0265_ clknet_leaf_68_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6005__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7817_ _1292_ _1296_ _3177_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8797_ _0196_ clknet_leaf_35_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7753__A1 _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7748_ _3110_ _3111_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_61_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _3018_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6308__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6492__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__I _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__C _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6244__A1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7744__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A2 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6369__C _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8666__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8472__A2 _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5286__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ _0381_ _0377_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6385__B _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4684__I _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8224__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6235__A1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5038__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ _1728_ _1415_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8720_ _0119_ clknet_leaf_50_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5932_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8651_ _0050_ clknet_leaf_35_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5863_ _0902_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7735__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6538__A2 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7602_ _2644_ _2969_ _2970_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__A1 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _4240_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8582_ _3864_ _3866_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5794_ _1327_ _3920_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7533_ as2650.pc\[6\] _0727_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _4245_ _4063_ _4221_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_108_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7464_ _1037_ as2650.stack\[5\]\[4\] as2650.stack\[4\]\[4\] _0942_ _2836_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4676_ _4255_ _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6415_ _1786_ _1799_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4859__I _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7395_ _2619_ _2766_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6710__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net52 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6346_ _1777_ _1802_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4721__A1 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6277_ as2650.stack\[2\]\[2\] _1746_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8016_ as2650.stack\[5\]\[9\] _3352_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5228_ _4048_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7671__C2 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__B _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5159_ _0551_ _0637_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7726__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8849_ _0248_ clknet_leaf_29_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6314__I _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5201__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7854__B _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8689__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8151__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__B1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7145__I _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4712__A1 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6984__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8454__A2 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4718__B _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7009__A3 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__A2 _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7965__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7965__B2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4779__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8390__A1 _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7193__A2 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7764__B _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6940__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4530_ _4021_ _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4461_ _4041_ _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6200_ _1121_ _1458_ _1693_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7180_ _2558_ _1635_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4392_ _3914_ _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6894__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _1624_ _0866_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8445__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5259__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ as2650.psl\[6\] _1539_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__B _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5013_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6208__A1 _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6964_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8703_ _0102_ clknet_leaf_33_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1439_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6895_ _2293_ _1274_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8634_ _0033_ clknet_leaf_3_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5846_ _1371_ _0660_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7184__A2 _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8831__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7674__B _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5195__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _1245_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8565_ _4202_ _2323_ _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6931__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__C _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7393__C _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7516_ as2650.stack\[2\]\[5\] _2792_ _0925_ as2650.stack\[3\]\[5\] _0975_ _2887_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4728_ _4285_ _4190_ _4156_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8496_ _2576_ _2425_ _3070_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8133__A1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7447_ _2031_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4659_ _4057_ _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6695__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7378_ _2653_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6329_ _0823_ _0829_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8436__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7849__B _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7947__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7568__C _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4856__S1 _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6044__I _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8372__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8372__B2 _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7584__B _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6979__I _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5883__I _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A3 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6922__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8124__A1 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8124__B2 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__I _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5110__A1 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8704__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__I _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_29_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__I _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8854__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__A2 as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5700_ _1234_ _1214_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ as2650.stack\[4\]\[2\] _2124_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7166__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8363__A1 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7494__B _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ as2650.stack\[5\]\[6\] _1165_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5793__I _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6913__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5716__A3 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8350_ _1189_ _1540_ _3643_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4924__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _1081_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _4205_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4513_ _4079_ _4092_ _4093_ _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8281_ _2904_ _3590_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5493_ _0687_ _0990_ _0991_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7232_ _2604_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7874__B1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4444_ as2650.ins_reg\[2\] _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7163_ _2267_ _2356_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4375_ _3912_ _3955_ _3927_ _3929_ _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__8418__A2 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6114_ _1104_ _1593_ _1608_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_101_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7094_ _2469_ _2478_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__B2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5033__I _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7929__A1 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7929__B2 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7996_ as2650.stack\[6\]\[1\] _1231_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6601__A1 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7157__A2 as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8354__A1 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _1327_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8617_ _0016_ clknet_leaf_27_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _1157_ _1339_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6904__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__A1 _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8548_ _1717_ _3795_ _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8479_ _3757_ _3767_ _3771_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8727__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7880__A3 _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5891__A2 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7093__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6039__I _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6840__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8877__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7396__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7148__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8345__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4906__A1 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7489__B _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4692__I _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7850_ _1387_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7387__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__A1 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6801_ as2650.r123\[3\]\[5\] _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5398__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7781_ _2265_ _2462_ _2723_ _3137_ _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4993_ _4226_ _0552_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5398__B2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6732_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7936__C _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8336__A1 _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7139__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ _1910_ _2111_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8402_ _3541_ _3698_ _3706_ _3296_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ _1126_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _2006_ _2021_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7952__B _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _3987_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8333_ _3391_ _3635_ _3640_ _3441_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8264_ _0730_ _0725_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5476_ as2650.stack\[3\]\[12\] as2650.stack\[0\]\[12\] as2650.stack\[1\]\[12\] as2650.stack\[2\]\[12\]
+ _0929_ _0978_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6114__A3 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4427_ _4007_ _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4867__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5322__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7215_ _1575_ _2274_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8195_ _2323_ _3506_ _3507_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7243__I _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ _1734_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5873__A2 _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ _3938_ _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7077_ _2461_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6028_ _1293_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5698__I _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8575__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8575__B2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7979_ _1487_ _3325_ _3330_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6050__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8327__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8327__B2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6889__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7550__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7838__B1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__A2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5864__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7066__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6992__I _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6813__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8566__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_80 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_91 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _4043_ _0883_ _0887_ _4277_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _0790_ _0793_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7000_ _1556_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5192_ _0747_ _0749_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7998__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7057__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7902_ _3242_ _3259_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6280__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5311__I _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8882_ _0281_ clknet_leaf_41_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7833_ _3192_ _3193_ _1257_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7764_ _2817_ _3078_ _2867_ _3053_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8309__A1 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _0331_ _0535_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7780__A2 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ as2650.stack\[3\]\[7\] _1754_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5791__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7695_ _2741_ _3060_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7238__I _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ as2650.r123_2\[2\]\[6\] _1948_ _2096_ _2043_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5543__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6577_ _0557_ _1995_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8316_ _3483_ _3622_ _3623_ _3624_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5528_ _1015_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8247_ _0658_ _3427_ _3550_ _3432_ _3557_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_59_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ _1012_ as2650.stack\[7\]\[11\] as2650.stack\[6\]\[11\] _1007_ _0954_ _1013_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8178_ _1663_ _0385_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7048__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ _1431_ _1099_ _2485_ _2512_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7599__A2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6271__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8548__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7220__A1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6023__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5782__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6052__I _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5534__A1 _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__S _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4888__A3 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7287__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A3 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4300__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7039__A1 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8539__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_2_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7211__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6014__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4830_ _0389_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7762__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4761_ _0323_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4576__A2 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _1954_ _1820_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7480_ _1160_ _2850_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4692_ _4271_ _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6431_ _0415_ _0788_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5525__A1 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _1818_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8101_ _2353_ _3415_ _3416_ _2609_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5313_ _4139_ _4140_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6293_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ _0781_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8032_ as2650.stack\[4\]\[9\] _3361_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _0562_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7450__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7450__B2 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8865_ _0264_ clknet_leaf_68_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7202__A1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ _1246_ _2598_ _2291_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8796_ _0195_ clknet_leaf_35_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5764__A1 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7747_ _3088_ _3056_ _1219_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4959_ _4166_ _0420_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7678_ _3043_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5516__A1 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _2015_ _2055_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__A2 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6047__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6244__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5886__I _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5755__A1 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__A1 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6180__B2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6235__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6980_ _1107_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__A2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _1184_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5796__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5994__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8172__I _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8650_ _0049_ clknet_leaf_35_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7735__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7601_ as2650.stack\[2\]\[7\] _1006_ _2797_ as2650.stack\[3\]\[7\] _2970_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4813_ _4237_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8581_ _1635_ _3865_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5793_ _1239_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _2610_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4744_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7499__A1 _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7463_ _2529_ _2823_ _2834_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4675_ _4254_ _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6414_ _0655_ _1210_ _1782_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8610__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7394_ _2620_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6345_ _1780_ _1801_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4721__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6276_ _1481_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8347__I _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7671__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8015_ _1113_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4875__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8760__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5158_ _0674_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7423__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5089_ _0552_ _0638_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__B _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8082__I _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8848_ _0247_ clknet_leaf_48_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8779_ _0178_ clknet_leaf_76_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__B2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7870__B _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4712__A2 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7662__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7414__A1 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__A2 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7965__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5728__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7193__A3 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7764__C _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8633__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__A1 _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6940__A3 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6240__I _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _3970_ _4040_ _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6153__A1 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _3909_ _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4703__A2 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5900__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6130_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__B1 _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _1381_ _1553_ _1554_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7071__I _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5012_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7405__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6208__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7956__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _2360_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8702_ _0101_ clknet_leaf_30_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ as2650.r123_2\[3\]\[0\] _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__C _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6894_ _1091_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8633_ _0032_ clknet_leaf_2_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5845_ _4025_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5195__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8564_ _2635_ _1406_ _2319_ _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5776_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7515_ _2788_ _2885_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4727_ _3940_ _4092_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8495_ _1717_ _3756_ _3772_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__I _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7446_ _1095_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6144__A1 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _4228_ _4230_ _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6695__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7892__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7377_ _2745_ _2747_ _2749_ _2750_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_104_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _4144_ _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _0789_ _0828_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7644__B2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ _1733_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8656__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4630__A1 _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7865__B _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8372__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7584__C _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7156__I _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6060__I _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8124__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6995__I _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7635__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4449__A1 _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5110__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7399__B1 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8363__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6374__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5561_ _1087_ _1092_ _1065_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7300_ _2313_ _1409_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ _4021_ _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8280_ _2855_ _2907_ _3528_ _2856_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5492_ _1036_ _0966_ _1043_ _1019_ _0983_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_144_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7874__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6677__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7231_ _2606_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7874__B2 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4443_ _4002_ _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4374_ as2650.cycle\[0\] _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7162_ _2484_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7015__B _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _0436_ _1379_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7093_ _2470_ _2476_ _2477_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5314__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6044_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8679__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__A1 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ _2116_ _3339_ _3340_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6946_ _1376_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6877_ _1288_ _1320_ _2277_ _1266_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_50_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7157__A3 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8354__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8616_ _0015_ clknet_leaf_60_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5828_ _1356_ _1340_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6365__A1 _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8547_ _3266_ _3834_ _3835_ _2279_ _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5759_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4915__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6117__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _2601_ _3768_ _3770_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7865__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__A2 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7429_ _2801_ _2758_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5891__A3 _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8290__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5643__A3 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4851__A1 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A1 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7595__B _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8345__A2 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6356__A1 _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5159__A2 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4906__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4303__I _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6659__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7856__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__C _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5331__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8821__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6831__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8033__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6800_ _2212_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8584__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7780_ _1272_ _2383_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5398__A2 as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _4234_ _0445_ _0421_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _0906_ _1827_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8336__A2 _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _0861_ _1910_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8401_ _1314_ _3702_ _3705_ _3588_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _1036_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _2025_ _2028_ _2023_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8332_ _3423_ _3639_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5544_ as2650.addr_buff\[7\] _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8263_ net34 _3572_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_133_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5475_ _0951_ as2650.stack\[7\]\[12\] as2650.stack\[6\]\[12\] _0920_ _0973_ _1028_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_117_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A4 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7214_ _1714_ _2234_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4426_ _3927_ _3932_ _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8194_ _2293_ _3488_ _2769_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7145_ _2527_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4357_ _3937_ _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _1090_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5086__A1 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _1518_ _1521_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7399__C _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8575__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6586__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7978_ as2650.stack\[7\]\[9\] _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _2319_ _2322_ _2324_ _2326_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6050__A3 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8090__I _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A1 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7862__C _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__A1 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7838__B2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__A1 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8844__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5864__A3 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8263__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7066__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5889__I _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6813__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8265__I _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A1 _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8566__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_70 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_81 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_92 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8318__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7829__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5260_ _0816_ _0801_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6501__A1 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5191_ _0747_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5855__A3 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8254__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7057__A2 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7901_ _1344_ _3240_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8881_ _0280_ clknet_leaf_40_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8557__A2 _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7832_ _1806_ _4118_ _2633_ _3990_ _1304_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_110_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7763_ _2502_ _3124_ _3125_ _2428_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4975_ _4156_ _0519_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8309__A2 _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8717__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6714_ _2136_ _1757_ _2148_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5791__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7694_ as2650.addr_buff\[2\] _2679_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7963__B _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6645_ _1899_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5543__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8867__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6576_ _2025_ _2028_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6740__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__B _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8315_ _2414_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _1071_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_121_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8246_ _2063_ _3456_ _3397_ _3556_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8493__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6099__A3 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _0950_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8493__B2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4409_ _3989_ _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8177_ _1954_ _0385_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7128_ _2408_ _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7048__A2 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5059__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7059_ _2447_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8548__A2 _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7756__C2 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7220__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5782__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7592__C _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6731__A1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5534__A2 _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4788__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8484__A1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8484__B2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7039__A2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5412__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__B _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8539__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6243__I _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4760_ _0321_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_61_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6970__A1 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5773__A2 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _4270_ _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _0824_ _1884_ _1885_ _1796_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6722__A1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6361_ _3890_ _4001_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_128_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7074__I _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8100_ _3221_ _2299_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5312_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8475__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6292_ _1753_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5289__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8031_ _2117_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5243_ _0782_ _0794_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7802__I _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8227__A1 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5174_ _0675_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8864_ _0263_ clknet_leaf_67_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7815_ _1069_ _1085_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7202__A2 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8795_ _0194_ clknet_leaf_36_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7746_ _1219_ _3088_ _3056_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6961__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5764__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7693__B _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7677_ _1204_ _1536_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4889_ _4075_ _0295_ _0383_ _0447_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_6628_ _2052_ _2054_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5516__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6174__C1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8301__C _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _2007_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4401__I _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8466__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8229_ _3242_ _3540_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7441__A2 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8154__B1 _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7108__B _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__I _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6012__B _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6180__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4311__I as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8209__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__A2 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7778__B _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5443__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ _1012_ _1078_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7196__A1 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7069__I _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7196__B2 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7600_ _0945_ as2650.stack\[1\]\[7\] as2650.stack\[0\]\[7\] _0942_ _2969_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4812_ _0374_ _4067_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8580_ _3790_ _2429_ _2430_ _3863_ _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5792_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6943__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _2897_ _2900_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4743_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__I _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7462_ _2828_ _2831_ _2833_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7499__A2 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4674_ as2650.r0\[2\] _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6413_ _1867_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7393_ _4010_ _2758_ _2765_ _2720_ _2392_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5317__I _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8448__A1 _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _1784_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8775__D _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6275_ _1134_ _1744_ _1745_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8014_ _3350_ _1193_ _3351_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5226_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5480__C _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7671__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _0650_ _0584_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5088_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8847_ _0246_ clknet_leaf_48_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6934__A1 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8778_ _0177_ clknet_leaf_76_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7729_ _1018_ _2977_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6611__I _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5227__I _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6162__A2 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7870__C _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7662__A2 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7178__A1 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4306__I _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8222__B _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6153__A2 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4390_ _3907_ _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5900__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7102__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7102__B2 _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input8_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5664__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ as2650.r123\[0\]\[5\] as2650.r123_2\[0\]\[5\] _3886_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7405__A2 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6962_ _2220_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7020__C _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8701_ _0100_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5913_ _1369_ _1424_ _1436_ _1438_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7169__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6893_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7169__B2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8632_ _0031_ clknet_leaf_2_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5844_ _1253_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6916__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8563_ _3754_ _2442_ _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5775_ _3909_ _3982_ _3973_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6392__A2 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ _2794_ as2650.stack\[1\]\[5\] as2650.stack\[0\]\[5\] _2789_ _2885_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4726_ _4297_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5475__C _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8494_ _3242_ _3785_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7445_ as2650.addr_buff\[4\] _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_120_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4657_ _3924_ _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6144__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7376_ _2648_ as2650.stack\[7\]\[2\] as2650.stack\[6\]\[2\] _0918_ _0971_ _2750_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4588_ _4167_ _4168_ _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6327_ _1782_ _1783_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5655__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5209_ _0766_ _0767_ _0626_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _1546_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6080__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4630__A2 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6907__A1 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4933__A3 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7332__A1 _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6135__A2 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7635__A2 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4449__A2 _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7399__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8217__B _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7399__B2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8060__A2 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__I _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5949__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5177__A3 _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6374__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8750__CLK clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7571__B2 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__I _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _4205_ _1100_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5295__C _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4511_ _4091_ _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7323__A1 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5491_ _1039_ _1040_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_144_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7323__B2 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7230_ _2605_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4442_ _3926_ _4014_ _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5885__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _3916_ _2356_ _1242_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7082__I _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4373_ _3953_ _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6112_ _1247_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7092_ _1402_ _2472_ _1593_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6043_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7994_ as2650.stack\[6\]\[0\] _1231_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _0495_ _2342_ _1606_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__A2 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6876_ _2271_ _2272_ _1319_ _2276_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7157__A4 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8615_ _0014_ clknet_leaf_58_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5827_ _0639_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7257__I _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7562__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__A2 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6161__I _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1260_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8546_ _3266_ _4251_ _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4471__S1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4709_ _4288_ _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7314__A1 _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8477_ _2361_ _1092_ _1262_ _3769_ _2594_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6117__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5689_ _1194_ _1224_ _1225_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7428_ _1594_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5325__B1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7865__A2 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__A2 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7359_ _2628_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5891__A4 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5628__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8623__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8042__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7876__B _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A2 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8773__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7595__C _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7553__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6356__A2 _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__A1 _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__A2 _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8502__B1 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4520__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7856__A2 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5619__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8281__A2 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4842__A2 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8033__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8584__A3 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4991_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _2152_ _2155_ _2162_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6661_ _2104_ _1858_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7077__I _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8400_ _3401_ _3704_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5612_ _1150_ _1155_ _1156_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6592_ _2003_ _2044_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8331_ _3636_ _3638_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5543_ _4154_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8262_ net51 _3545_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _0967_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5858__A1 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _2334_ _2350_ _2588_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4425_ _4005_ _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8193_ _3407_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8646__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7144_ _1255_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4356_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _2293_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8272__A2 _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6026_ _4280_ _0861_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8796__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4833__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8024__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7696__B _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6586__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7977_ _3326_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5995__I _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4597__A1 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _0436_ _1386_ _2325_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_126_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7535__A1 _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6859_ _3919_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6889__A3 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5010__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8529_ _4169_ _4182_ _0299_ _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6510__A2 _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4521__A1 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8566__A3 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_60 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A2 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_71 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_82 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_93 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_127_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8669__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7829__A2 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__A2 _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ as2650.holding_reg\[6\] _3940_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8254__A2 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7360__I _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5068__A2 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8006__A2 _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7900_ _3245_ _3255_ _3257_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8880_ _0279_ clknet_3_1_0_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6017__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7831_ _2216_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8405__B _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7765__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7765__B2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7762_ _2263_ _2462_ _2918_ _3123_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4974_ _0527_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5240__A2 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6713_ as2650.stack\[3\]\[6\] _1754_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7693_ _3056_ _3058_ _2501_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7517__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5791__A3 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7517__B2 _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6644_ _0769_ _2094_ _1817_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _1968_ _2026_ _2027_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8140__B _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6740__A2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8314_ net35 _3389_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5526_ _1073_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__B2 _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8245_ _3551_ _3554_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5457_ _1007_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6099__A4 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ as2650.ins_reg\[5\] _3945_ _3947_ _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8176_ _3401_ _3488_ _2484_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5388_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _3931_ _2235_ _2487_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__I _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _3918_ _3919_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8245__A2 _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7058_ _2446_ _0627_ _2421_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4806__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _1503_ _0738_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7756__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A2 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7756__B2 _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4990__A1 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8811__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8181__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6731__A2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8484__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8236__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6247__A1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8209__C _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7995__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4309__I _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6970__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _4269_ _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A3 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6360_ _3993_ _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4733__A1 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _4097_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6291_ _1754_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8475__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8030_ _1478_ _3359_ _3360_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5242_ _0795_ _0798_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4928__B _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8227__A2 _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ _4018_ _0716_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6789__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7986__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8932_ net46 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8863_ _0262_ clknet_leaf_66_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7738__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7814_ _1256_ _1273_ _2523_ _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_8794_ _0193_ clknet_3_6_0_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8834__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7745_ _2261_ _3078_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4957_ _4189_ _0420_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6961__A2 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8163__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ as2650.pc\[10\] _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4888_ _0378_ _4231_ _0369_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_123_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _0870_ _2050_ _2011_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6174__B1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6174__C2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6713__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6558_ _0666_ _1233_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5509_ _0870_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6489_ _1919_ _1943_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8466__A2 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8228_ net32 _3483_ _3539_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8096__I _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8159_ _3444_ _2713_ _2714_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7729__A1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5204__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6952__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4963__A1 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8154__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8154__B2 _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7901__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8457__A2 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7903__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8707__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8209__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6640__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _3991_ _1378_ _0910_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _1308_ _1317_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6943__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7530_ _1170_ _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4954__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4742_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8402__C _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7461_ _2784_ _2832_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4673_ _4080_ _4252_ _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6412_ _1777_ _1802_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4706__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _2761_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6343_ _1786_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8448__A2 _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6274_ as2650.stack\[2\]\[1\] _1498_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5225_ as2650.r123\[0\]\[6\] as2650.r123_2\[0\]\[6\] as2650.psl\[4\] _0784_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8013_ as2650.stack\[5\]\[8\] _1165_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5156_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7969__B _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8791__D _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _0626_ _0630_ _0644_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8846_ _0245_ clknet_leaf_48_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8384__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8777_ _0176_ clknet_leaf_77_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6934__A2 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _1207_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7728_ _3074_ _3091_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4945__A1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8136__B2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8312__C _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__B _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7659_ _3001_ _3003_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6698__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7723__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__I _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8127__A1 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8222__C _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__A3 _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4322__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7102__A2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6249__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _3883_ _0569_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_85_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6861__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5664__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6613__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6961_ _2356_ _2358_ net26 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8700_ _0099_ clknet_leaf_46_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5912_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6892_ _1283_ _1309_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8366__A1 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8366__B2 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8631_ _0030_ clknet_leaf_23_wb_clk_i as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ as2650.psu\[5\] _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6916__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7808__I _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8562_ _3230_ _3845_ _3847_ _3849_ _2493_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5774_ _1248_ _1266_ _1279_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_7513_ _2533_ _2875_ _2883_ _2743_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4725_ _4162_ _0288_ _4137_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5328__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8493_ _0978_ _3780_ _3784_ _3772_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7444_ _2313_ _1591_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4656_ _4232_ _4235_ _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5352__A1 _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _4139_ _4140_ _3938_ _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7375_ _2644_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ _0580_ _0831_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6257_ _1416_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _0753_ _0676_ _0489_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5655__A2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7699__B _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6188_ _1646_ _1682_ _0439_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5139_ _0414_ _0304_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__C _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7211__C _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6080__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8829_ _0228_ clknet_leaf_28_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6907__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8109__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7580__A2 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A3 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5343__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6540__B1 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5894__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7402__B _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7399__A2 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4317__I _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4385__A2 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4510_ _4084_ _4090_ _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _0976_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8520__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _4021_ _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4987__I _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7160_ _2539_ _2541_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_78_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5885__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4372_ _3935_ _3936_ _3952_ _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7087__A1 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6111_ _1069_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _2471_ _2272_ _2472_ _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6834__A1 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6042_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8127__C _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8587__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7993_ _3338_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6062__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6944_ _2314_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8339__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6875_ _1247_ _1421_ _2238_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__8143__B _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8614_ _0013_ clknet_leaf_58_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5826_ _1349_ _1353_ _1355_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8545_ _3789_ _1624_ _3833_ _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5757_ _3934_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ _4286_ _4287_ _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8476_ _1402_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7314__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8511__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ as2650.stack\[6\]\[12\] _1202_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7427_ _2653_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5325__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _4219_ _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5876__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7358_ _2397_ _2727_ _2731_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7078__A1 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ as2650.stack\[3\]\[14\] _1765_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7289_ _2660_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6825__A1 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8578__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__A1 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7876__C _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7002__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7553__A2 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7305__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8502__A1 _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5867__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6816__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5619__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7241__A1 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4990_ _4228_ _0420_ _0445_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6660_ _0886_ _1900_ _1857_ _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_108_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6347__A3 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ as2650.stack\[5\]\[4\] _1135_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5555__A1 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _1949_ _2029_ _2042_ _2043_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8330_ _3637_ _3612_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5542_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8261_ _3390_ _3570_ _3571_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5473_ _0943_ as2650.stack\[5\]\[12\] as2650.stack\[4\]\[12\] _0968_ _1026_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5606__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7212_ _2584_ _2587_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4424_ _4004_ _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5858__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8192_ _1396_ _2945_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7143_ _1244_ _1425_ _2525_ _2470_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4355_ _3896_ _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7074_ _2375_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7480__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6025_ _0647_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5341__I _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7976_ _1478_ _3325_ _3328_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7783__A2 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5794__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__A2 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _4009_ _1588_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7268__I _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6858_ _1660_ _2246_ _2262_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5809_ _0442_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__A4 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _2114_ _2191_ _2195_ as2650.r123_2\[1\]\[7\] _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6900__I _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A3 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _4169_ _4182_ _0300_ _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7299__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8459_ _2470_ _1727_ _3753_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8248__B1 _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A2 _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__B1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7471__A1 _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7887__B _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6026__A2 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_61 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_72 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_83 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A1 _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6015__C _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6810__I _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4760__A2 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__I _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6501__A3 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7641__I _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7214__A1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6017__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7830_ _1093_ _3920_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8557__A4 _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7761_ _1227_ _3110_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _0532_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4505__I _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6712_ _2133_ _1757_ _2147_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7692_ _3042_ _3057_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _0722_ _1951_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5528__A1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8613__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ _1971_ _1988_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8313_ _2994_ _3421_ _3616_ _3452_ _3621_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xclkbuf_leaf_22_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5525_ _4174_ _0575_ _0911_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4751__A2 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8244_ _3551_ _3554_ _3189_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ _1009_ as2650.stack\[5\]\[11\] as2650.stack\[4\]\[11\] _0946_ _1010_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6876__B _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8794__D _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4407_ _3901_ _3987_ _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8175_ net31 _3487_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5700__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ _0922_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _2507_ _2509_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4338_ as2650.addr_buff\[5\] _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7453__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7057_ _2063_ _2376_ _1426_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6008_ _0856_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6008__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7756__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7959_ _3311_ _3248_ _3312_ _0904_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__I _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7508__A2 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7692__A1 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7444__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6077__I _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7995__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8225__C _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8636__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8879__D _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4981__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6183__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7380__B1 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8786__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__I _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5310_ _0736_ _0549_ _0864_ _4233_ _0867_ _4128_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_142_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6290_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6486__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4995__I _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5241_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A1 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5172_ _4264_ _0551_ _0637_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8227__A3 _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7435__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5446__B1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7986__A2 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_8931_ net47 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8416__B _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8862_ _0261_ clknet_leaf_15_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7813_ _1270_ _1594_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A1 _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8793_ _0192_ clknet_leaf_36_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7744_ _3009_ _3107_ _2954_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _0516_ _4166_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8151__B _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7675_ _1198_ _2849_ _3041_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7546__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4887_ _0446_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6626_ _2048_ _2055_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6174__A1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6174__B2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6557_ _2008_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5066__I _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5508_ as2650.r123\[0\]\[7\] _0963_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6488_ _1922_ _1942_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8227_ _3480_ _3534_ _3538_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7674__A1 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_1_1_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5439_ as2650.stack\[3\]\[10\] _0934_ _0937_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8158_ net30 _3471_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6229__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _2414_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8089_ _1395_ _2945_ _2301_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5988__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8659__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7729__A2 _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4412__A1 _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4963__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7901__A2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7665__A1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7191__I _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__B2 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__B1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6640__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _4256_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _3975_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4741_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4954__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7460_ _2031_ _2227_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7353__B1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _4081_ _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _1780_ _1801_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4706__A2 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7391_ _2715_ _2717_ _2763_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6342_ _1791_ _1795_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7656__A1 _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _1484_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8012_ _1122_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5224_ _4085_ _0573_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _0668_ _0670_ _0672_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8801__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5086_ _0489_ _0645_ _0317_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8146__B _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8845_ _0244_ clknet_leaf_48_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8384__A2 _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8776_ _0175_ clknet_leaf_76_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7592__B1 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _1487_ _1483_ _1489_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7727_ _2946_ _3083_ _3073_ _2667_ _1414_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_40_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4945__A2 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4939_ _0403_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6147__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7658_ _2852_ _3024_ _2954_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6609_ _1831_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6698__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7589_ _2956_ _2929_ _2957_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_1_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_88_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4881__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6355__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5189__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7886__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7638__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__I _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8824__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6861__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4872__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8063__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6265__I _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _1327_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4624__A1 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _4187_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6891_ _3946_ _2289_ _2290_ _1438_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8366__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8630_ _0029_ clknet_leaf_27_wb_clk_i as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5842_ _1349_ _1367_ _1368_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6377__A1 _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8561_ _3848_ _3830_ _1688_ _1502_ _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5773_ _1290_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7096__I _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7512_ _1427_ _2876_ _2628_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4724_ _4138_ _4139_ _4140_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6129__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8492_ _2528_ _0927_ _3783_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7443_ _1152_ _2773_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4655_ _4233_ _4227_ _4234_ _4231_ _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_116_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7374_ _2645_ as2650.stack\[5\]\[2\] as2650.stack\[4\]\[2\] _1008_ _2748_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _4138_ _4166_ _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7629__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6325_ _0796_ _0821_ _1781_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6256_ _1105_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5104__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6884__B _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _0753_ _0287_ _0676_ _0765_ _0344_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_76_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7699__C _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6187_ _1680_ _1681_ _1429_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _4049_ _0573_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ as2650.holding_reg\[5\] _0584_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4615__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6903__I _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6368__A1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8828_ _0227_ clknet_leaf_26_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7565__B1 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8759_ _0158_ clknet_leaf_1_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4918__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8109__A2 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4423__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7317__B1 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7868__A1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8847__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8045__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6085__I _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__A2 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8348__A2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7909__I _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7020__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5031__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7859__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8520__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4440_ _4015_ _3898_ _3965_ _4020_ _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5334__A2 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _3941_ _3951_ _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6110_ _1072_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8284__A1 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7087__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _1377_ _1382_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6834__A2 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6041_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6196__S _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8036__A1 as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8587__A2 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7992_ _1185_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _1298_ _2222_ _1609_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8424__B _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6723__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _2273_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8613_ _0012_ clknet_leaf_58_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5825_ net45 _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__A4 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8544_ _4214_ _2354_ _3832_ _1530_ _1561_ _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5756_ _1281_ _4186_ _1284_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_72_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4707_ _4165_ _4084_ _4090_ _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8475_ _1411_ _1579_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5687_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7426_ _2791_ _2793_ _2796_ _2798_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_135_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4638_ _4218_ _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6522__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7357_ _2728_ _2730_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4569_ _4100_ _4046_ _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7078__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8275__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _1497_ _1763_ _1766_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7288_ _2662_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6825__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6239_ _1530_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8027__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8578__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4418__I _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5636__I0 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__A2 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__A3 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__I _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7002__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6761__A1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__A2 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6816__A2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8018__A1 as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7132__C _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8569__A2 _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__B _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5004__A1 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ _1828_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5555__A2 _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__I _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5541_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ net51 _3418_ _3321_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ _0557_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6504__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5307__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7211_ _1611_ _2585_ _2586_ _1608_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4423_ as2650.ins_reg\[3\] _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8191_ _3489_ _3500_ _3503_ _3443_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5858__A3 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8257__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7142_ _2522_ _2524_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4354_ _3926_ _3934_ _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7073_ _2455_ _2457_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8009__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _0348_ _0491_ _0547_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__7480__A2 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7975_ as2650.stack\[7\]\[8\] _3327_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6926_ _2323_ _0896_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6991__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5794__A2 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8692__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6857_ _2261_ _2253_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5808_ _1328_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6788_ _2205_ _2206_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6743__A1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8527_ _3815_ _0492_ _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5739_ _3960_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6402__B _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7284__I _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7299__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8496__A1 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8458_ _2258_ _1726_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7409_ _2391_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8389_ net38 _3654_ _3655_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8248__A1 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8248__B2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5532__I _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7471__A2 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7887__C _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4592__B _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8064__B _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5234__A1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_62 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_73 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_84 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5785__A2 _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5537__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5707__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8487__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8239__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__B2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__A2 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7369__I _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6273__I _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7760_ _1227_ _3098_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _0284_ _0332_ _0469_ _0323_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6973__A1 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6711_ as2650.stack\[3\]\[5\] _2143_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7691_ _1198_ _3029_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6642_ _2036_ _2091_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6725__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5528__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _1971_ _1988_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8312_ _2389_ _3619_ _3620_ _2952_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8478__A1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5524_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8243_ _3514_ _3552_ _3515_ _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_5455_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4406_ _3982_ _3986_ _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_62_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8174_ net30 net29 net28 _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5386_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8149__B _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7125_ _2288_ _2475_ _2508_ _2235_ _3931_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4337_ as2650.addr_buff\[6\] _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7453__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _2445_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6007_ _4174_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8402__A1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__B _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7958_ _1636_ _3248_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6909_ _3900_ _3997_ _4076_ _4267_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7889_ _1528_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7508__A3 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__A2 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__C1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7913__B1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4990__A3 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7141__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4587__B _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6358__I _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7444__A2 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5207__B2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4606__I _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7917__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A2 _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7380__A1 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5437__I _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7380__B2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7132__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7652__I _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__S _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _0665_ _4218_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4497__B _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6268__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _0729_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5446__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8930_ net47 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_110_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8416__C _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8861_ _0260_ clknet_leaf_18_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4516__I _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7812_ _0898_ _2316_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8792_ _0191_ clknet_3_6_0_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _2902_ _3100_ _3106_ _2504_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4955_ as2650.holding_reg\[4\] _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7674_ _2896_ _3039_ _3040_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4886_ _0383_ _4234_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8151__C _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6625_ _2045_ _2057_ _2075_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6174__A2 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8730__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4804__S0 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _1975_ _1976_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5507_ _1057_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7123__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6487_ _1926_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8226_ _2857_ _3416_ _3537_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8880__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5685__A1 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8157_ net52 net28 _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5369_ _0921_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _2458_ _2491_ _2492_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8088_ _3391_ _3399_ _3403_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _4293_ _2422_ _2431_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6937__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A2 _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8568__I _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7665__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4479__A2 _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5428__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8517__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5720__I _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8603__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8753__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4740_ as2650.r123\[0\]\[1\] as2650.r123_2\[0\]\[1\] _3886_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4671_ _4075_ _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7353__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5167__I _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7353__B2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6410_ _1773_ _1864_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7390_ _2762_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6341_ _1793_ _1796_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7105__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _1121_ _1495_ _1743_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8011_ _2138_ _3345_ _3349_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5667__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5223_ _0698_ _0702_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ _4035_ _0687_ _0713_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5419__A1 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6726__I _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5085_ as2650.holding_reg\[5\] _0584_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6092__A1 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6919__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8844_ _0243_ clknet_leaf_49_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8162__B _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7592__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8775_ _0174_ clknet_3_2_0_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5987_ as2650.stack\[2\]\[9\] _1488_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7726_ _2362_ _3079_ _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4938_ _0373_ _0307_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7657_ _2902_ _3017_ _3023_ _2504_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6147__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _0337_ _4263_ _4229_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ as2650.r123_2\[2\]\[5\] _1830_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7588_ net3 _4101_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7895__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _0422_ _1903_ _1843_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8209_ _0424_ _0453_ _3466_ _3490_ _3491_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8626__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4330__A1 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7241__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6083__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5830__A1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8776__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7895__C _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7583__A1 _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6138__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7886__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5897__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5715__I _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6310__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7151__B _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8063__A2 _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7810__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A2 _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _1425_ _1435_ _1424_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6890_ net22 _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ net21 _1354_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6377__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ _1293_ _1297_ _1298_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8560_ _0861_ _1514_ _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7511_ _2879_ _2881_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4723_ _4192_ _4171_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8491_ _3781_ _3782_ _2528_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6129__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7442_ _2619_ _2813_ _2767_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7877__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4654_ _4228_ _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7373_ as2650.stack\[2\]\[2\] _1006_ _0926_ _2746_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_122_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4585_ _4165_ _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5625__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__A3 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6324_ _0666_ _0306_ _0822_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8649__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7629__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4560__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6255_ _1730_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6301__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _0473_ _0749_ _0757_ _0325_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6186_ _1636_ _1301_ _1418_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4685__B _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8799__CLK clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7061__B _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5137_ _0619_ _0695_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8054__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__B1 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _0627_ _0585_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4615__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8827_ _0226_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8758_ _0157_ clknet_leaf_1_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _2618_ _3073_ _2777_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7317__B2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8689_ _0088_ clknet_leaf_43_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8514__B1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5423__S0 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8293__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7750__I _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8067__B _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6366__I _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8045__A2 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5803__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5031__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A1 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7925__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5319__B1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7859__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4370_ _3943_ _3950_ _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6040_ net2 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__A3 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8036__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7795__A1 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7991_ _1500_ _3333_ _3337_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6942_ _1317_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_16_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ _3949_ _1250_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8612_ _0011_ clknet_leaf_58_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5824_ _1325_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5755_ _4122_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8543_ _2323_ _3790_ _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4706_ _4285_ _4188_ _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5686_ _0615_ _1211_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8474_ _3758_ _3760_ _3761_ _3766_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8511__A3 _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] _3887_ _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7425_ as2650.stack\[2\]\[3\] _0918_ _2797_ as2650.stack\[3\]\[3\] _0975_ _2798_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__6522__A2 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7356_ _1138_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4568_ _4103_ _4052_ _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6307_ as2650.stack\[3\]\[13\] _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7287_ _1129_ _1116_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _4044_ _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6286__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _1715_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8027__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ as2650.psl\[7\] _1299_ _1663_ as2650.overflow _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6038__A1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7786__A1 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6589__A2 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5636__I1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6914__I _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A4 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4434__I _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6210__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8350__B _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8266__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6277__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4609__I _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8018__A2 _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7226__B1 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7529__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4344__I _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5004__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8260__B _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _1088_ _3986_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4763__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5471_ as2650.r123\[0\]\[4\] _0987_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5307__A3 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7701__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _1612_ _2326_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4422_ _4002_ _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8190_ _2761_ _3502_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ _1573_ _2523_ _2518_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8257__A2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4353_ _3933_ _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5903__I _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7072_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7323__C _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _4183_ _0301_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4519__I _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7768__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6734__I _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _3326_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5243__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8837__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__S1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6925_ _1645_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ as2650.addr_buff\[4\] _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ _1328_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8170__B _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _0806_ _1949_ _2195_ as2650.r123_2\[1\]\[6\] _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7940__A1 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8601__D _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8526_ _0462_ _0850_ _3814_ _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5738_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8457_ _0496_ _2103_ _3752_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8496__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5669_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7408_ _2778_ _2739_ _2779_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8388_ _3042_ _3422_ _3693_ _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8396__I _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8248__A2 _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7339_ as2650.pc\[1\] net6 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5813__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7208__B1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output45_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A1 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A2 _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A3 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_63 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_74 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_85 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4993__A1 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7931__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__A1 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__B _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6498__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6819__I _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8239__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__I _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__C _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5473__A2 as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4971_ _0475_ _0472_ _0529_ _0530_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_63_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6973__A2 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _2130_ _2141_ _2146_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8175__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7690_ _1205_ _1197_ _3029_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_32_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _0726_ _2036_ _1836_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7922__A1 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6725__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4802__I _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _2023_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8311_ _2994_ _3566_ _2660_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5523_ _4007_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7686__B1 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5454_ _0941_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8242_ _1674_ _0555_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4405_ _3983_ _3985_ _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__A1 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8173_ _3420_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5385_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5633__I _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4336_ _3907_ _3916_ _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7124_ _1425_ _1401_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7989__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _2444_ _0516_ _2421_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6661__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _0845_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_31_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8402__A2 _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7957_ as2650.psu\[7\] _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4975__A1 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6908_ _0638_ _0661_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7888_ _1533_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7509__B _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6839_ _2244_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6177__B1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5808__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7913__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__C2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7913__B2 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A1 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8509_ _0473_ _4279_ _3798_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8469__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7141__A2 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7898__C _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5207__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7601__B1 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A3 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6707__A2 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7132__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5453__I _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__A1 _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5170_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__8682__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6643__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_65_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8860_ _0259_ clknet_leaf_16_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7811_ _1717_ _1529_ _3157_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8791_ _0190_ clknet_leaf_0_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7742_ _2614_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4957__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _4225_ _0493_ _0515_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6159__B1 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7673_ _2581_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4885_ _0428_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6624_ _2046_ _2056_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7371__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4804__S1 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _1935_ _2007_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5506_ _1047_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7123__A2 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6486_ _1929_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8225_ _1152_ _3405_ _3536_ _2720_ _2660_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5437_ _0374_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5363__I _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8156_ _2404_ _3469_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5368_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ _1437_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ _3899_ _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8087_ _3400_ _3402_ _2484_ _2612_ _1318_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5299_ _0856_ _4107_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6634__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7038_ _1600_ _2419_ _2429_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_56_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8139__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8139__B2 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5538__I _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7898__B1 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7362__A2 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8311__A1 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5273__I _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8517__C _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8378__A1 _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6928__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7050__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__B _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ _4093_ _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7353__A2 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8550__A1 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6340_ _4254_ _0786_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8302__A1 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6271_ as2650.stack\[2\]\[0\] _1498_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6864__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5222_ _0703_ _0709_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8010_ as2650.stack\[6\]\[7\] _3338_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7612__B _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5153_ as2650.r123\[1\]\[5\] _0600_ _0712_ _0408_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__I _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6616__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _0344_ _0629_ _0643_ _4148_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_110_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6092__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8843_ _0242_ clknet_leaf_26_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6919__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8774_ _0173_ clknet_leaf_77_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1484_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7592__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7725_ _2345_ _3087_ _3089_ _2916_ _2467_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ _0497_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _2945_ _3022_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4868_ _4262_ _4260_ _4265_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8541__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _1949_ _2058_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5355__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7587_ _2083_ _0669_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _3888_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6538_ _0433_ _1821_ _1991_ _1956_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6189__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7647__A3 _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _4096_ _0831_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8208_ _0424_ _0453_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4330__A2 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8139_ _2669_ _3422_ _3451_ _3453_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_114_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5821__I _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6607__A1 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6083__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5594__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8599__B2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7151__C _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7271__A1 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8720__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7023__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ _4107_ _1329_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8870__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _1301_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5178__I _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ _2391_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _4299_ _0284_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8490_ _2695_ _1593_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8523__A1 _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7441_ _2611_ _2807_ _2812_ _2302_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4653_ _4127_ _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4810__I _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ as2650.stack\[1\]\[2\] as2650.stack\[0\]\[2\] _0928_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4584_ _4025_ _4004_ _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5127__B _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6323_ _0819_ _1778_ _1779_ _0830_ _0838_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_131_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _1725_ _1727_ _1716_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5205_ _4157_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6185_ _1418_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _0417_ _4220_ _0502_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7262__A1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__B2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ as2650.holding_reg\[5\] _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5812__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7014__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8826_ _0225_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6368__A3 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__A2 _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8757_ _0156_ clknet_leaf_1_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5576__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5088__I _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _1224_ _1473_ _1474_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7708_ _3072_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8688_ _0087_ clknet_leaf_43_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8514__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8514__B2 _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7639_ _2801_ _2991_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5879__A2 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__S1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4551__A2 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8743__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5500__B2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6056__A2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7478__I _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6382__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5111__S0 _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8505__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__A1 _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__B2 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5726__I _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8102__I _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7941__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6834__A4 _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5461__I _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7990_ as2650.stack\[7\]\[14\] _3335_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7795__A2 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _2336_ _2338_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _1645_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8611_ _0010_ clknet_leaf_58_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5823_ _1350_ _1339_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6755__B1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8542_ _1571_ _3830_ _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5754_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8616__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7337__B _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4705_ as2650.holding_reg\[1\] _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8473_ _1392_ _2368_ _3763_ _3765_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5685_ _1221_ _1214_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4540__I _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7424_ _0925_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4636_ _4199_ _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8766__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7355_ _1130_ _2673_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5730__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ _4028_ _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ _1756_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7286_ _2660_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8168__B _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4498_ _4031_ _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7483__A1 _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6237_ _1310_ _1714_ _1081_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5371__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6168_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6038__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5119_ _0655_ _4247_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6099_ _4122_ _1376_ _1594_ _1374_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5797__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5549__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8809_ _0208_ clknet_leaf_64_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6210__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5546__I _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7474__A1 _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6277__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7474__B2 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7226__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7226__B2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7777__A2 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5788__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7001__I _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8639__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7529__A2 _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4763__A2 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8789__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4360__I _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _1004_ _1023_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6996__B _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _4001_ _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5712__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7140_ _1373_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4352_ _3927_ _3932_ _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7465__A1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ _3955_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6022_ _0769_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7217__A1 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7768__A2 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7973_ _3323_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4535__I _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6924_ _2226_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5243__A3 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6991__A3 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6855_ _2260_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5806_ _1326_ _1337_ _1338_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6786_ _2096_ _2197_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7940__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8525_ _0850_ _1345_ _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5737_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8456_ _0890_ _3734_ _3736_ as2650.r123\[2\]\[7\] _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5668_ _0501_ _1158_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ _2778_ _2739_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4619_ _3999_ _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8387_ _3679_ _3692_ _2400_ _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5599_ _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7338_ _2710_ _2711_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5315__B _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7269_ _0944_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7208__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6925__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7208__B2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4445__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_53 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_75 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_86 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_26_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6195__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6195__B2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A2 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5942__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7695__A1 _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__A1 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__I _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4970_ _0322_ _0468_ _0477_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_75_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _1048_ _1839_ _2088_ _2090_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6186__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6571_ _2004_ _2005_ _2022_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_121_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8310_ _2994_ _2297_ _3562_ _3618_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5522_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7686__A1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8241_ _1674_ _0555_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7686__B2 _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5453_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4404_ as2650.cycle\[3\] _3984_ _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8172_ _3480_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7334__C _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5384_ _0935_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7123_ _2377_ _2372_ _2503_ _2506_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4335_ _3915_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7989__A2 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8804__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7054_ _1660_ _2441_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6005_ _1500_ _1495_ _1501_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6661__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71_wb_clk_i clknet_opt_1_1_wb_clk_i clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7956_ _3260_ _0862_ _3308_ _3309_ _1525_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_36_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6907_ _3931_ _2304_ _2305_ _1635_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7576__I _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7887_ _3207_ _0492_ _3226_ _3244_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6838_ as2650.addr_buff\[0\] _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6177__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__B2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7913__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5096__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _1861_ _2191_ _2193_ as2650.r123_2\[1\]\[0\] _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8508_ _1247_ _2591_ _1420_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8439_ _3735_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5824__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7429__A1 _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6101__A1 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7260__B _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6404__A2 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5207__A3 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7486__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8157__A2 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A4 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7904__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7668__A1 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7668__B2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5734__I _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__I _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7154__C _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6340__A1 _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8827__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__A1 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__I _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6643__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7840__A1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 io_in[5] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7810_ _3158_ _1335_ _3170_ _1550_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8790_ _0189_ clknet_leaf_36_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4406__A1 _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _3103_ _3104_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ as2650.r123\[1\]\[3\] _4212_ _0514_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4957__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7672_ _3017_ _3025_ _3038_ _2982_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6159__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4884_ _4229_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6159__B2 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6623_ _2061_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5906__A1 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _0580_ _1792_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4969__B _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7659__A1 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5505_ _0771_ _0990_ _0991_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6485_ _1930_ _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8320__A2 _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8224_ _2777_ _2811_ _3506_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _0962_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6331__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8155_ _3465_ _3468_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5367_ _0922_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7106_ _2459_ _2480_ _2490_ _1421_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4318_ as2650.ins_reg\[4\] _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8086_ _3401_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8176__B _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5298_ as2650.holding_reg\[7\] _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _0310_ _2397_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7831__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7939_ _3152_ _0726_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5819__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8139__A2 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7347__B1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7898__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7898__B2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5554__I _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8311__A2 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5125__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6873__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4884__A1 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7702__C _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8378__A2 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7050__A2 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5729__I _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4633__I _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__C _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8550__A2 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7105__A3 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6270_ _1742_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5221_ _0704_ _0778_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8066__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5152_ _0690_ _0693_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7813__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6616__A2 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5083_ _0331_ _0634_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4627__A1 _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6092__A3 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8842_ _0241_ clknet_leaf_27_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8773_ _0172_ clknet_leaf_76_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _1200_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7724_ _3088_ _3056_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4936_ _0400_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ _3018_ _3021_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _0428_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8541__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6606_ _2045_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7586_ _2852_ _2953_ _2954_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5355__A2 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _0353_ _0354_ _0355_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6537_ _0426_ _1821_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _1210_ _1882_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8207_ _0561_ _3456_ _3397_ _3518_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5419_ _0936_ _0933_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_79_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ _4062_ _1835_ _1837_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8057__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8138_ _3452_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6607__A2 _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7804__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8069_ _3383_ _3384_ _1429_ _2229_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_43_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7032__A2 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8672__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8800__D _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6543__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5897__A3 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6846__A2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__B2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8048__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8220__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7023__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4363__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _1302_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6782__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _4291_ _4175_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7440_ _2614_ _2811_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4652_ _4127_ _4227_ _4229_ _4231_ _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7371_ as2650.stack\[3\]\[2\] _0934_ _0937_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _4016_ _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _0823_ _0829_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8287__B2 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6253_ _1728_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8039__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5204_ _0752_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6184_ _1636_ _1647_ _1648_ _1659_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _0618_ _0620_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7262__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _0317_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8695__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__A1 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8825_ _0224_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6773__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8756_ _0155_ clknet_leaf_43_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5576__A2 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ as2650.stack\[1\]\[12\] _1469_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ _1213_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _0470_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8687_ _0086_ clknet_leaf_30_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5899_ _1370_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8514__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7638_ _2743_ _3005_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6525__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5879__A3 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7569_ _2934_ _2935_ _2937_ _2938_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6828__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__I _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8450__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__A3 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8364__B _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8202__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__C _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5111__S1 _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__A1 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7308__A3 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4911__I _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8505__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5742__I _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4358__I _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6940_ _1647_ _1581_ _2337_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_66_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6871_ _1274_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5007__A1 _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8610_ _0009_ clknet_leaf_59_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5822_ _1351_ _1340_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6755__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5753_ _1285_ _1286_ _1097_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7618__B _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8541_ _0862_ _1514_ _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4704_ _4143_ _4145_ _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6507__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8472_ _2466_ _3764_ _2328_ _3131_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5684_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7423_ _2788_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4635_ _4215_ _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7180__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7354_ _2501_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _4146_ _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5730__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6305_ _1494_ _1763_ _1764_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7285_ _1278_ _1611_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _4070_ _4072_ _4074_ _4077_ _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6236_ _1300_ _1408_ _1713_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7483__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6167_ _0351_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8432__A1 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5118_ _4022_ _0422_ _0664_ _0677_ _3954_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6038__A3 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _1263_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5049_ _0365_ _0305_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8808_ _0207_ clknet_leaf_66_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5549__A2 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8739_ _0138_ clknet_leaf_58_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5827__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7171__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8710__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7171__B2 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7710__A3 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7263__B _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7226__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__A1 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8423__B2 _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5237__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5511__B _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6393__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7631__C1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6985__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5788__A2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4460__A2 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6737__A1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5737__I _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6061__C _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4420_ _3999_ _4000_ _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_126_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5712__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4351_ _3929_ _3931_ _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5472__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7070_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4523__I0 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _1516_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8414__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7217__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6976__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7972_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _4194_ _1398_ _1399_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_35_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _2258_ _2259_ _2245_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout49 net13 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5805_ net42 _1333_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7348__B _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6785_ _2203_ _2204_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ _1072_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8524_ _0747_ _1518_ _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5951__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7153__A1 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8455_ _0496_ _2082_ _3732_ _0771_ _3751_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5667_ _1205_ _1161_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7406_ _0423_ _0362_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4618_ _4198_ _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8386_ _2544_ _3682_ _3691_ _3281_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ as2650.pc\[3\] _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5703__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8179__B _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7083__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7337_ _1130_ _1118_ _1139_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4549_ _4055_ _4129_ _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7268_ _2643_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7811__B _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6219_ _1466_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7199_ _1432_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8405__A1 _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7208__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_54 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_26_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_65 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A1 _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8361__C _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__I _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4745__A3 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5942__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7772__I _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7695__A2 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8089__B _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7447__A2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8606__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4636__I _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8108__I _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7012__I _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8552__B _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8756__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__B _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7383__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _2004_ _2005_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5521_ _1069_ net10 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _0657_ _0654_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5146__B1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5452_ _0921_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7686__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ as2650.cycle\[2\] _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8171_ _3482_ _3484_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5383_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7122_ _2504_ _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4334_ _3909_ _3911_ _3914_ _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_99_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7053_ _1350_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6110__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6004_ as2650.stack\[2\]\[14\] _1498_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__B _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6949__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7610__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7955_ _3205_ _0868_ _3207_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ net23 _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7886_ _2564_ _0460_ _3243_ _2547_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6837_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6177__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_40_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8507_ _1320_ _1582_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7126__A1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5719_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6699_ as2650.stack\[3\]\[0\] _1765_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7677__A2 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8438_ _3738_ _1897_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5688__A1 as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8369_ net50 _3636_ _3638_ _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7429__A2 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8629__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6101__A2 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8779__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5860__A1 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4456__I _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7601__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6340__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A1 _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8093__A2 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5750__I _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5851__A1 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4366__I as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 io_in[6] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_83_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__B _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4406__A2 _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7740_ as2650.pc\[12\] _2083_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4952_ _0496_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7671_ _0981_ _2752_ _3024_ _3037_ _3031_ _2623_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_4883_ _0318_ _0319_ _0363_ _0368_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_60_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6159__A2 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _2059_ _2060_ _2073_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5906__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5462__S0 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _1979_ _1981_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8305__B1 _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5504_ _1048_ _0914_ _1054_ _1019_ _0958_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_69_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4590__A1 _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7659__A2 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6484_ _1934_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8223_ _1269_ _3532_ _2819_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5435_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6331__A2 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A1 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ as2650.psu\[1\] _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8154_ _1532_ _3192_ _3467_ _3922_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4893__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7105_ _1614_ _2488_ _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4317_ _3897_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8085_ _3911_ _1294_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ _0325_ _0847_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7036_ _1531_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7831__A2 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A4 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _3292_ _3293_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7347__A1 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7869_ _3152_ _0386_ _3227_ _2547_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8544__B1 _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7898__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4879__C _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4333__A1 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4884__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6086__A1 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__A1 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5011__S _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4850__S _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8121__I _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4572__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7510__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _0581_ _4221_ _0707_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5151_ _0694_ _0697_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8066__A2 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7813__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5082_ _0482_ _0636_ _0641_ _0287_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4627__A2 _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8841_ _0240_ clknet_leaf_22_wb_clk_i as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8772_ _0171_ clknet_leaf_76_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1478_ _1483_ _1486_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7723_ as2650.pc\[11\] _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4935_ as2650.r0\[1\] _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7654_ _3019_ _2988_ _3020_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _0363_ _0368_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ _2046_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7585_ _2620_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4797_ _0354_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6536_ _1771_ _1989_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7501__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6467_ _1876_ _1920_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6304__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8206_ _3456_ _3517_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5418_ _0951_ as2650.stack\[7\]\[9\] as2650.stack\[6\]\[9\] _0920_ _0973_ _0974_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_6398_ _1840_ _1854_ _1835_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4866__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8137_ _2287_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5349_ _4000_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8057__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5323__C _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8068_ _1241_ _2818_ _1249_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5815__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7019_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7568__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7568__B2 _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8817__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7740__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8296__A2 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6396__I _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4857__A2 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__I _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8048__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6854__I0 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8544__C _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _4295_ _4298_ _4297_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4793__A1 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _4230_ _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7731__A1 _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7370_ _2533_ _2732_ _2742_ _2743_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4582_ _4162_ _4142_ _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ _0823_ _0829_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6298__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6252_ _1416_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5203_ _0631_ _0632_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8039__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6183_ _1649_ _1671_ _1672_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5134_ _0617_ _0621_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5065_ _4225_ _0599_ _0625_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6470__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4554__I _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8824_ _0223_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8211__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8755_ _0154_ clknet_leaf_71_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5967_ _1464_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6773__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7970__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7706_ _1205_ _3014_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4784__A1 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4918_ _0346_ _0478_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8686_ _0085_ clknet_leaf_31_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5898_ _1384_ _1393_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7637_ _2498_ _3000_ _3004_ _2733_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7722__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4849_ _3888_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5385__I _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7722__B2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7568_ _0949_ as2650.stack\[7\]\[6\] as2650.stack\[6\]\[6\] _2792_ _0971_ _2938_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6519_ _1888_ _1972_ _1936_ _1937_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7499_ _2853_ _2857_ _2773_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6289__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__A3 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8450__A2 _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__A4 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5264__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6461__A1 _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__B1 _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8202__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8380__B _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7961__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6612__C _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8505__A3 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7713__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__A3 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8269__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4639__I _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A2 _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__A1 _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _2270_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ _0422_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7952__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8540_ _3813_ _3827_ _3828_ _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5752_ _3982_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4703_ _4126_ _4236_ _4278_ _4282_ _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8471_ _4164_ _4194_ _1102_ _1101_ _1254_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__7704__A1 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6507__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7422_ _2794_ as2650.stack\[1\]\[3\] as2650.stack\[0\]\[3\] _2789_ _2795_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4634_ _4214_ _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7180__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ _2723_ _2712_ _2718_ _2724_ _2726_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5191__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _4143_ _4145_ _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5933__I _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6304_ as2650.stack\[3\]\[12\] _1759_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7353__C _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4496_ _3967_ _4076_ _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7284_ _2606_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6235_ _1371_ _1085_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_65_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8662__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ as2650.psl\[3\] _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _4079_ _0676_ _4093_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6038__A4 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6097_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _4255_ _0498_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__A1 _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__B2 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8807_ _0206_ clknet_leaf_64_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7809__B _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6999_ _2366_ _2282_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7943__A1 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8738_ _0137_ clknet_leaf_44_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8669_ _0068_ clknet_leaf_24_wb_clk_i as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6939__I _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__I as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8120__A1 _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8806__D _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__A2 _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5237__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7631__C2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6985__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8187__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6849__I as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__A1 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4350_ _3930_ as2650.cycle\[0\] _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_125_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8685__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4920__A1 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8111__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _1509_ _1512_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4523__I1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6425__A1 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7971_ _3323_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ _1251_ _1401_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8178__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ as2650.addr_buff\[3\] _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4739__A1 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5804_ _0965_ _1329_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6784_ _0712_ _2188_ _2193_ as2650.r123_2\[1\]\[5\] _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8523_ _3794_ _3810_ _3812_ _3624_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5735_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8454_ as2650.r123\[2\]\[6\] _3736_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5666_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8350__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ _0352_ _4252_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4617_ _3935_ _4197_ _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8385_ _2404_ _3689_ _3690_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5597_ _1115_ _1142_ _1143_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__C _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7336_ _1137_ _1128_ as2650.pc\[0\] _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _4127_ _4128_ _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7267_ _2642_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _4057_ _4059_ _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5467__A2 _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6664__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _1121_ _1473_ _1703_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7198_ _2574_ _2575_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8405__A2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _1527_ _1547_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A2 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_55 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_88 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7916__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4742__I _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A4 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8341__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__B1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6655__A1 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6618__B _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A1 _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7168__C _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8580__A1 _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__A3 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ as2650.halted _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7135__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8332__A1 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__A1 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__B2 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _0410_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4402_ _3912_ as2650.cycle\[0\] _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5697__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8170_ net30 _3483_ _3224_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5382_ _0921_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7121_ _2229_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4333_ _3912_ _3913_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7052_ _2424_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _1236_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8399__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6949__A2 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8700__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7954_ _3153_ _0886_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6905_ _1421_ _2296_ _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7885_ _2569_ _0454_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6836_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8571__A1 _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8850__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _1769_ _2190_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _1428_ _3795_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5718_ _1082_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6698_ _2138_ _2131_ _2139_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8437_ _4185_ _3733_ _3737_ _3739_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5393__I _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8368_ _3485_ _3673_ _3674_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8087__B1 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ _2505_ _2693_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8299_ _0875_ _2104_ _3607_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_105_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6637__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7541__C _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7113__I _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5860__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5568__I _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8562__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8562__B2 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5376__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8314__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4351__A2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8547__C _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8723__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput7 io_in[7] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_65_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7053__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__B1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5603__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4951_ _0509_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4382__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7670_ _2743_ _3036_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4882_ _0410_ _4066_ _0441_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ _2061_ _2043_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7907__B _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5462__S1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6552_ _1923_ _1987_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8305__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8305__B2 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5119__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5503_ _1050_ _1051_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6483_ _1936_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4590__A2 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8222_ _3525_ _3533_ _2300_ _3226_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6867__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5434_ _0908_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6331__A3 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7642__B _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4342__A2 _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8153_ _2255_ _0386_ _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5365_ as2650.psu\[0\] _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6619__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7104_ _1728_ _2342_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4316_ _3890_ _3896_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8084_ net28 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5296_ _4157_ _0849_ _0853_ _4027_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7292__A1 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7035_ _1272_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7044__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7595__A2 _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7937_ _1157_ _3240_ _3224_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7868_ _3152_ _0393_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7347__A2 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8544__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8544__B2 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6819_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7799_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6858__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__I _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8746__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4333__A2 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5530__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4467__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__A2 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7283__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8383__B _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6682__I _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6615__C _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__A1 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8535__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4930__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4572__A2 _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7018__I _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7510__A2 _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8558__B _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _0703_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8066__A3 _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__I _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5081_ _0336_ _0639_ _0640_ _4176_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8471__B1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4627__A3 _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7026__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8840_ _0239_ clknet_leaf_24_wb_clk_i as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8771_ _0170_ clknet_leaf_78_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5983_ as2650.stack\[2\]\[8\] _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7722_ _2816_ _3083_ _3072_ _2379_ _3086_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_75_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ _4023_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8619__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5001__I _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7653_ _1188_ _1537_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4865_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ _2049_ _2055_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _2611_ _2944_ _2952_ _2302_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4796_ _0338_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8769__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6535_ _1968_ _1971_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_88_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _1879_ _1892_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8468__B _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8205_ _1660_ _0556_ _3516_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_122_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__A1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6397_ _1842_ _1844_ _1852_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8136_ _3442_ _3446_ _3450_ _1571_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ _0894_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8067_ _2223_ _2237_ _2312_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5279_ _0835_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5276__B1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _4187_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7017__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6776__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6007__I _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8517__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7547__B _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4750__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6170__C _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7740__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8378__B _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5581__I _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5806__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6854__I1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__I _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7559__A2 _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6231__A2 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8508__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _4047_ _4053_ _4083_ _4089_ _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput10 wb_rst_i net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4581_ _4161_ _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6320_ _0832_ _0837_ _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7495__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6251_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5202_ _0629_ _0759_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6182_ _0425_ _0523_ _1649_ _4201_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _0608_ _0691_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5064_ as2650.r123\[1\]\[4\] _0600_ _0624_ _0408_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6470__A2 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8823_ _0222_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8211__A3 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8754_ _0153_ clknet_leaf_55_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5966_ _1217_ _1465_ _1472_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7705_ _2271_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4917_ _0284_ _0332_ _0324_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8685_ _0084_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5897_ _1396_ _1403_ _1411_ _1422_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_139_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7636_ _3001_ _3003_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _0366_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7722__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__A2 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7567_ _2643_ _2936_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7881__I _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _0331_ _0334_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _0416_ _1792_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _2723_ _2851_ _2861_ _2724_ _2868_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _0872_ _1844_ _1902_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__A4 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8119_ _4068_ _4130_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7121__I _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__B2 _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__B1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6764__A3 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7961__A2 _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7713__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5724__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7791__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7477__A1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5820_ _0557_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8290__C _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7952__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ as2650.cycle\[3\] _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4281_ _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8470_ _1419_ _3762_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5682_ as2650.pc\[12\] _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7421_ _0922_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4633_ _4063_ _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7352_ _2256_ _2634_ _2725_ _2281_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _3997_ _4144_ _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7468__A1 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _1754_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7283_ _1119_ _2607_ _2658_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4495_ _4017_ _4075_ _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5479__B1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6234_ _1179_ _1467_ _1712_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8807__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6691__A2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6165_ _1655_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _3957_ _1251_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7640__A1 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _0604_ _0606_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4454__A1 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__A2 _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8806_ _0205_ clknet_3_1_0_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7809__C _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6998_ _1258_ _2272_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7097__B _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8737_ _0136_ clknet_leaf_58_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5949_ as2650.stack\[0\]\[13\] _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8668_ _0067_ clknet_leaf_24_wb_clk_i as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7619_ _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8599_ as2650.psu\[3\] _3878_ _3880_ _3870_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8500__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7459__A1 _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__A2 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6131__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6955__I _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4693__A1 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7631__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6985__A3 _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8187__A2 _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7934__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4920__A2 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6122__A1 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6673__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6865__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7217__A4 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7622__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7970_ _1112_ _1183_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4436__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6976__A3 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ _3902_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8178__A2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _1533_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5803_ _1335_ _1330_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6783_ _2061_ _2072_ _2197_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8522_ as2650.psl\[5\] _3811_ _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5734_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7689__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8453_ _0687_ _3732_ _3749_ _3750_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5665_ as2650.pc\[10\] _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8350__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _2229_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _4196_ _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8384_ _1295_ _3676_ _2407_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5164__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6361__A1 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ as2650.stack\[5\]\[2\] _1135_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7335_ _2605_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4547_ _3976_ as2650.idx_ctrl\[0\] _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_89_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7266_ _0917_ _0924_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6113__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _4058_ _3919_ _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_1_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6664__A2 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ as2650.stack\[1\]\[0\] _1475_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7197_ _2538_ _1240_ _1633_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _1101_ _1250_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7613__A1 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _4005_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_56 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7916__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__I _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8230__I _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6352__A1 _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6104__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__B2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8386__B _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6685__I _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7852__A1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7604__A1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7080__A2 _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7907__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8580__A2 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6591__A1 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8652__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8332__A2 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ as2650.r123\[0\]\[3\] _0963_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6343__A1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4401_ _3929_ _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5381_ as2650.stack\[3\]\[8\] _0934_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7120_ _2301_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4332_ as2650.cycle\[0\] _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_114_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6646__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7843__A1 _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7051_ _2424_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _1497_ _1495_ _1499_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6949__A3 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7953_ _3203_ _3306_ _3307_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5082__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6904_ _2297_ _1276_ _2292_ _2298_ _2300_ _2302_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8315__I _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7884_ _1437_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6835_ _2225_ _2232_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5909__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ _2190_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6582__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5717_ _3900_ _4145_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8505_ _1570_ _1431_ _2473_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5674__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ as2650.stack\[4\]\[7\] _2134_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8323__A2 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5648_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8436_ _3738_ _1804_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6334__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6885__A2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8367_ net50 _3654_ _3655_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8087__A1 _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7318_ _2617_ _2663_ _2692_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8087__B2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8298_ _3605_ _3582_ _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7834__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _2344_ _2466_ _2499_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7834__B2 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__A3 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5849__I _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4753__I _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8675__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8562__A2 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6325__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7522__B1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6876__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8078__A1 _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7732__C _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7825__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7304__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5300__A2 _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 io_in[8] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8250__A1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__A2 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5759__I _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4950_ _0510_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8002__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4881_ _4250_ _0442_ _4247_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6620_ _2062_ _1833_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_33_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6551_ _1982_ _1986_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8305__A2 _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5502_ _0977_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6316__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _0579_ _0788_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8221_ _2408_ _3528_ _3529_ _3532_ _3423_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6867__A2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ as2650.r123\[0\]\[2\] _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4878__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6331__A4 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8152_ _2250_ _4242_ _4243_ _3428_ _3429_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_5364_ _0917_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7103_ _2482_ _2485_ _2487_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6619__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4315_ _3895_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8083_ _2564_ _3393_ _3395_ _3398_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5295_ _0850_ _0737_ _0852_ _0473_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7034_ _4138_ _2422_ _2427_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7292__A2 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8698__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8241__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__A2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5055__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__I _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7936_ _2306_ _3198_ _3282_ _3291_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7867_ _1293_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8544__A2 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6818_ _1095_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6555__A1 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__B1 _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7798_ _1563_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6749_ _2157_ _1031_ _2160_ _1025_ _2166_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7833__B _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8419_ _3425_ _3721_ _3722_ _3391_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7552__C _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7807__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8480__A1 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__A3 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6963__I _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8232__A1 _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__I _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7794__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8535__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7727__C _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6546__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__A3 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7743__B _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5521__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6078__C _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5080_ _0627_ _0336_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8840__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8471__A1 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8471__B2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5285__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8574__B _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8223__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7026__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8770_ _0169_ clknet_leaf_78_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5588__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7721_ _1410_ _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7918__B _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4933_ _4143_ _0494_ _4194_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_33_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8526__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7652_ _2983_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6537__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4864_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _2052_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7583_ _2946_ _2951_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _0356_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_59_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6534_ _1923_ _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _1879_ _1892_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8204_ _3514_ _3515_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5416_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6396_ _1807_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5512__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8135_ _2669_ _3406_ _3449_ _3412_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5347_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8066_ _2159_ _2592_ _3380_ _3381_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__8462__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5278_ as2650.r0\[7\] _4219_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5276__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7017_ _2263_ _2400_ _2412_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5276__B2 _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8214__A1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7017__A2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5028__A1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7919_ _1351_ _3221_ _3273_ _3275_ _3202_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8517__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8713__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6958__I _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7055__S _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8863__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6700__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8205__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8508__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7029__I _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ as2650.psl\[3\] as2650.carry _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8569__B _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6250_ _4037_ _1612_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7495__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _0645_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4388__I _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6181_ _1673_ _0871_ _0675_ _0729_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8444__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5132_ _0603_ _0622_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _0601_ _0602_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_84_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4856__I1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8822_ _0221_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5012__I _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8753_ _0152_ clknet_leaf_55_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5965_ as2650.stack\[1\]\[11\] _1469_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8736__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7704_ _2453_ _3069_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4916_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8684_ _0083_ clknet_leaf_25_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5896_ _1414_ _1375_ _1419_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_33_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7635_ _3002_ _2958_ _1095_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7183__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ _4225_ _0396_ _0409_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _0287_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7566_ _2794_ as2650.stack\[5\]\[6\] as2650.stack\[4\]\[6\] _0941_ _2936_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6930__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6517_ _1919_ _1969_ _1970_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5682__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ _2217_ _2866_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _0442_ _1903_ _1843_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ _4119_ _4124_ _1819_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8118_ _3189_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5249__A1 _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8049_ _3323_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6997__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8199__B1 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6749__B2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__C _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__B2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8609__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8426__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8759__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4671__I _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5750_ _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _3926_ _4279_ _4280_ _3992_ _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_72_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5681_ _1187_ _1217_ _1218_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4632_ as2650.r123\[1\]\[0\] _4212_ _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7420_ _0949_ as2650.stack\[7\]\[3\] as2650.stack\[6\]\[3\] _2792_ _0971_ _2793_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6912__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _2255_ _1268_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4563_ _3947_ _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _1492_ _1755_ _1762_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7282_ _2608_ _2657_ _2582_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4494_ _4054_ _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5479__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6233_ as2650.stack\[1\]\[7\] _1464_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8417__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1650_ _1658_ _1648_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6095_ _1311_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5046_ _0605_ _0507_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7640__A2 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4454__A2 _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5651__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8805_ _0204_ clknet_leaf_67_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6997_ _1327_ _2393_ _1100_ _4279_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4581__I _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_74_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__C _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8736_ _0135_ clknet_leaf_59_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5948_ _1451_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8667_ _0066_ clknet_leaf_35_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _1102_ _4027_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_90_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7618_ _2943_ as2650.pc\[6\] _1536_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8598_ _3879_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7549_ _2265_ _2818_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7459__A2 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8408__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A2 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4756__I _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7631__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6971__I _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7395__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8592__B1 _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__I _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A1 _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6658__B1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7751__B _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6122__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__I3 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5881__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__I _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8138__I _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A2 as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6881__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6976__A4 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6920_ _2316_ _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _2255_ _2246_ _2257_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7386__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5497__I _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _0350_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _2201_ _2202_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5936__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8521_ _3796_ _3809_ _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5733_ _1094_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8452_ as2650.r123\[2\]\[5\] _3736_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5664_ _1187_ _1201_ _1203_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6897__B1 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7403_ _2354_ _2772_ _2775_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4615_ _4191_ _4195_ _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8383_ _2256_ _3687_ _3688_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5595_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6361__A2 _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4372__A1 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4546_ as2650.idx_ctrl\[1\] _3977_ _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7334_ _1130_ _2659_ _2708_ _2415_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7310__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ as2650.addr_buff\[6\] _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7265_ _2624_ _2625_ _2640_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6113__A2 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5960__I _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6216_ _1179_ _1452_ _1702_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7196_ _4010_ _2515_ _2571_ _2573_ _2454_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _1059_ _1626_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7613__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _1391_ _1406_ _1407_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _0377_ _0552_ _0553_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_57 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_79 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8719_ _0118_ clknet_leaf_49_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7129__A1 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5155__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6352__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__I _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8386__C _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7852__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6187__B _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__I _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7080__A3 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7368__A1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6591__A2 _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _3954_ _3968_ _3980_ _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4354__A1 _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8577__B _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ as2650.cycle\[1\] _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _2422_ _2439_ _2440_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7843__A2 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ as2650.stack\[2\]\[13\] _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7952_ _1167_ _3197_ _3040_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7883_ _3239_ _3241_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _2233_ _1323_ _2234_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__8020__A2 _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5020__I _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6765_ _4202_ _1827_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6582__A2 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__I _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8504_ _2280_ _3793_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5716_ _4025_ _4120_ _4192_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6696_ _1178_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5176__B _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8435_ _4199_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5647_ as2650.pc\[8\] _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A1 _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8366_ _3028_ _3486_ _3668_ _3453_ _3672_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7317_ _2625_ _2674_ _2691_ _1430_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8087__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4529_ _4095_ _4107_ _4109_ _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8297_ _1538_ _0721_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6098__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7248_ _2609_ _1729_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7834__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__A2 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7179_ _1302_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7598__A1 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7770__A1 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__I _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7058__S _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5086__B _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6325__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7522__B2 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6876__A3 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8078__A2 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7825__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5836__A1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput9 io_in[9] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8250__A2 _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7320__I _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5064__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8538__B1 _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8002__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4880_ _0338_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6013__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7476__B _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ as2650.r123_2\[2\]\[4\] _1830_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5772__B1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5501_ as2650.stack\[3\]\[14\] as2650.stack\[0\]\[14\] as2650.stack\[1\]\[14\] as2650.stack\[2\]\[14\]
+ _1014_ _1015_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7513__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _1931_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4327__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8220_ net32 _3531_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5432_ _0962_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8069__A2 _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8151_ _1532_ _3456_ _3398_ _3464_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5363_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _2268_ _2486_ _3950_ _3916_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _3894_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7816__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8082_ _3397_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5294_ as2650.holding_reg\[7\] _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ _2423_ _2426_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4854__I _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8241__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7230__I _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__A2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7935_ _1356_ _3221_ _3202_ _3290_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7866_ _3223_ _3225_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6817_ _1073_ _1107_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7752__A1 _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6555__A2 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7797_ _1566_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7752__B2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _2000_ _2164_ _2177_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7504__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6679_ _1141_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6307__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8418_ _2558_ _3718_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A2 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8349_ _3390_ _3653_ _3656_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8480__A2 _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8642__CLK clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7140__I _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7991__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8792__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7743__A1 _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5595__I _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8299__A2 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7743__C _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4939__I _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5809__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8471__A2 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6482__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4674__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8223__A2 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _1481_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7720_ _2783_ _3084_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _3896_ _3941_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4796__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7651_ as2650.pc\[9\] _0728_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__A2 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6602_ _2051_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4548__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5745__B1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7582_ _2947_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4794_ _4264_ _4234_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _1982_ _1986_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7934__B _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__B1 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _1874_ _1875_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8203_ _2824_ _0459_ _3459_ _3460_ _3494_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__4849__I _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5415_ _0952_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6170__B1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _0350_ _1812_ _1845_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_86_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8134_ _3132_ _2671_ _3408_ _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8665__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5346_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8065_ _2241_ _2322_ _2341_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8462__A2 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5277_ _0609_ _0833_ _0834_ _0791_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5276__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7016_ _2340_ _2406_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8214__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7422__B1 as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7918_ _1535_ _3247_ _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ _3150_ _0301_ _3155_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7725__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6528__A2 _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7725__B2 _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6700__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A2 _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6907__C _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5267__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A1 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4494__I _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8205__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6923__B _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6767__A2 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7964__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4778__A1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7716__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7754__B _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8688__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8141__A1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7045__I _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5200_ as2650.holding_reg\[5\] _0471_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _4269_ _0295_ _0421_ _1674_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _0603_ _0622_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8444__A2 _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5258__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6455__A1 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ _0603_ _0608_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_69_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6207__A1 as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8821_ _0220_ clknet_leaf_26_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_2_1_wb_clk_i_I clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7955__A1 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8752_ _0151_ clknet_leaf_54_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _1208_ _1465_ _1471_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7703_ _3042_ _2608_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5430__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4915_ _3938_ _0337_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8683_ _0082_ clknet_leaf_50_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5895_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7707__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7634_ _0874_ _4101_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4846_ as2650.r123\[1\]\[2\] _4212_ _0407_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7183__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8380__A1 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ as2650.stack\[2\]\[6\] _2792_ _2797_ as2650.stack\[3\]\[6\] _0975_ _2935_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _0336_ _0338_ _0339_ _4176_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6930__A2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6516_ _1922_ _1942_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8132__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7496_ _2263_ _2818_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6447_ _1811_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8495__B _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8117_ _3431_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5329_ _4114_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5249__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6446__A1 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8048_ _2123_ _3369_ _3370_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6997__A2 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8199__A1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8199__B2 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7946__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__I _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8371__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8830__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6969__I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4932__A1 _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8123__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__I _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8426__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6637__C _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5660__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7937__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4471__I0 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _3990_ _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ as2650.stack\[6\]\[11\] _1202_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8362__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4631_ _4211_ _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6879__I _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5176__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7570__C1 _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7350_ _2676_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4562_ _4026_ _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ as2650.stack\[3\]\[11\] _1759_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7281_ _2609_ _2622_ _2655_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4493_ _4073_ _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6232_ _1173_ _1467_ _1711_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8417__A2 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6163_ _1651_ _0425_ _1654_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7625__B1 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _1587_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8703__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _0605_ _0507_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5023__I _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5651__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7928__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4862__I _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8804_ _0203_ clknet_leaf_35_wb_clk_i as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _2391_ _1087_ _2392_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8853__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8735_ _0134_ clknet_leaf_58_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5947_ _1224_ _1458_ _1459_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8666_ _0065_ clknet_leaf_33_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8353__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ _4204_ _4005_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7617_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _0390_ _0380_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8597_ _1005_ _2355_ _3774_ _3246_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4914__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7548_ _2675_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8105__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7479_ _1151_ _1144_ _2710_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_134_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6131__A3 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8408__A2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6029__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7919__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__I _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7395__A2 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8592__B2 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8344__A1 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4905__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6370__A3 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6658__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6122__A3 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8726__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5881__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7083__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8280__B1 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8876__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__A3 as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6850_ _2256_ _2253_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7386__A2 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _1326_ _1332_ _1334_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6781_ _0624_ _2188_ _2193_ as2650.r123_2\[1\]\[4\] _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7993__I _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8520_ _2459_ _0548_ _3796_ _3809_ _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5732_ _1249_ _1259_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7926__C _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8335__A1 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8451_ _4217_ _2058_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5663_ as2650.stack\[6\]\[9\] _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8103__B _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6897__A1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ _2773_ _2774_ _2728_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4614_ _4192_ _4194_ _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8382_ _1296_ _3075_ _3686_ _3684_ _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5594_ _0993_ _1127_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7333_ _2661_ _2663_ _2707_ _2606_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4545_ _4125_ _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4372__A2 _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7264_ _2627_ _2628_ _2629_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _3918_ _4056_ _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7310__A2 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6215_ as2650.stack\[0\]\[7\] _1449_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8329__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5321__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _1240_ _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7233__I _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__A2 _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _1548_ _1626_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4507__S0 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6077_ _1410_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6821__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _0557_ _4247_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_58 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8574__A1 _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ _2273_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8718_ _0117_ clknet_leaf_26_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7129__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8326__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8649_ _0048_ clknet_leaf_32_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6888__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__A1 _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6812__A1 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5598__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7368__A2 _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8565__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7540__A2 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4354__A2 _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ as2650.cycle\[6\] _3910_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6000_ _1484_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7951_ _0733_ _1721_ _3297_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6902_ _1255_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7882_ _0993_ _3240_ _3224_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8556__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _2237_ _2238_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__B _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _4216_ _4223_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8308__A1 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8503_ _3266_ _3792_ _3288_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5715_ _1084_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5790__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6695_ _2136_ _2131_ _2137_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8434_ as2650.r123\[2\]\[0\] _3736_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5646_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8365_ _1736_ _3670_ _3671_ _3023_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4345__A2 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5577_ _1067_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8487__C _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7316_ _2361_ _2677_ _2683_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ as2650.psl\[3\] _4108_ _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8296_ _1538_ _0721_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7295__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6098__A2 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7247_ _2270_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4459_ _3906_ _3922_ _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7178_ _2453_ _2557_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7047__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _1257_ _0898_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6751__B _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7770__A2 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__I _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A2 _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5836__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7038__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8538__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7210__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6013__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7761__A2 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__B2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5500_ _1012_ as2650.stack\[7\]\[14\] as2650.stack\[6\]\[14\] _0940_ _0954_ _1051_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_119_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6480_ as2650.r0\[4\] _0784_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6887__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5431_ _0964_ _0986_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4327__A2 as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8150_ _3459_ _3462_ _3463_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5362_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _1321_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _3893_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8081_ _3396_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7816__A3 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5293_ _0335_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7032_ _1673_ _2398_ _2425_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6127__I _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ _1428_ _3247_ _3274_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7865_ _0965_ _3203_ _3224_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6004__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _1249_ _2218_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7796_ _1258_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6747_ as2650.r123_2\[0\]\[3\] _2165_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _2123_ _2119_ _2125_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8417_ _1297_ _3718_ _3719_ _3720_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5629_ _1167_ _1158_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5515__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__A3 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8348_ _3636_ _3654_ _3655_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8279_ _3423_ _3573_ _3587_ _3588_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5818__A2 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7440__A1 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6037__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7991__A2 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8252__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7743__A2 _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8456__B1 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7431__A1 _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7431__B2 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5980_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8590__C _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__B1 as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7982__A2 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _0457_ _0461_ _0492_ _4039_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_46_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4796__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__I _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7650_ _3014_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4862_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7734__A2 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ _4097_ _1233_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5745__A1 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7581_ _2948_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4548__A2 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5745__B2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _4092_ _4265_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _1984_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7498__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7498__B2 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6463_ _1870_ _1894_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8202_ _2824_ _0459_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5414_ _0967_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6170__A1 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ _4070_ _1847_ _1848_ _1849_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8133_ _2680_ _3447_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4720__A2 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8064_ _2653_ _2312_ _2317_ _3379_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _0415_ _0498_ _0613_ _4254_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7015_ _1570_ _2408_ _2368_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4865__I _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_68_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7670__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7422__A1 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7422__B2 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _1258_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5984__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8072__I _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ _2570_ _4236_ _3206_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7779_ as2650.pc\[14\] _3139_ _3140_ _2502_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7489__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7416__I _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__A2 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4775__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6195__C _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7413__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6216__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7964__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7100__B _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7716__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7770__B _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5130_ _0601_ _0688_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5290__B _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _0617_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4466__A1 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4856__I3 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8820_ _0219_ clknet_leaf_26_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7955__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8751_ _0150_ clknet_leaf_55_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4769__A2 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5966__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5963_ as2650.stack\[1\]\[10\] _1469_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7702_ _2982_ _3066_ _3067_ _3051_ _2605_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5430__A3 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ as2650.holding_reg\[2\] _3938_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7168__B1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5894_ _1280_ _1309_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8682_ _0081_ clknet_leaf_25_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7633_ as2650.addr_buff\[0\] _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4845_ _4199_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5718__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ _2788_ _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8632__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ as2650.holding_reg\[2\] _0335_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6391__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _1943_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7495_ _0658_ _2461_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__C _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _4267_ _1847_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6694__A2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7891__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8782__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ _3923_ _1819_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8116_ _1321_ _3191_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5328_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__I _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8047_ as2650.stack\[7\]\[1\] _3335_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5259_ _0782_ _0794_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4457__A1 _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8199__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5501__S0 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8371__A2 _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5185__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__A2 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7146__I _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6134__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7882__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4696__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7634__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6988__A3 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7937__A2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8655__CLK clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4471__I1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _4187_ _4199_ _4210_ _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5176__A2 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7570__C2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _4137_ _4141_ _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8114__A2 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6300_ _1490_ _1755_ _1761_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7280_ _2495_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4492_ _4023_ _4024_ _4030_ _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8596__B _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6231_ as2650.stack\[1\]\[6\] _1464_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7873__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4687__A1 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ as2650.psu\[4\] _1655_ _0729_ net27 _0915_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_124_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5113_ _0668_ _0670_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _1383_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5304__I _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5044_ _4245_ _4063_ _0307_ _0501_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8762__D _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8803_ _0202_ clknet_leaf_20_wb_clk_i as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6995_ _2370_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8734_ _0133_ clknet_leaf_59_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5946_ as2650.stack\[0\]\[12\] _1454_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8665_ _0064_ clknet_leaf_32_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5877_ _0538_ _1402_ _1370_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _2903_ _2947_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4828_ _4129_ _0383_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8596_ _2258_ _2441_ _3869_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7547_ _2914_ _2915_ _2916_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4759_ _0320_ _0318_ _0319_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4914__A2 _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8105__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6116__A1 _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7478_ _2606_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6429_ _1793_ _1797_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4678__A1 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4678__B2 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6419__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8678__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7919__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8041__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__I _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8592__A2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5884__I _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5158__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4905__A2 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7855__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7607__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A2 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8435__I _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A1 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ net41 _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6780_ _2042_ _2197_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ _1261_ _1262_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8450_ _0599_ _3732_ _3747_ _3748_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6346__A1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5662_ _1186_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7401_ _1137_ _2729_ _2757_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4613_ _4193_ _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6897__A2 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8381_ _3683_ _3684_ _3685_ _3686_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _1139_ _1131_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7332_ _2664_ _2706_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7942__C _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4544_ _3898_ _4119_ _4124_ _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4372__A3 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7263_ _2631_ _2636_ _1430_ _2638_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7846__A1 _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4475_ as2650.addr_buff\[5\] _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ _1173_ _1452_ _1701_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7194_ _2558_ _2561_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6145_ _4280_ _1639_ _1522_ _1516_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8820__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6076_ _1529_ _1545_ _1569_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4507__S1 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6821__A2 _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _4022_ _0523_ _0566_ _0587_ _4065_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A1 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_59 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6585__A1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ _1687_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8717_ _0116_ clknet_leaf_25_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _1446_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7129__A3 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8080__I _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8648_ _0047_ clknet_opt_3_0_wb_clk_i as2650.r123_2\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6888__A2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8579_ as2650.psl\[1\] _3863_ _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4899__A1 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7852__C _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8262__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7065__A2 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5076__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8014__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__A3 _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8565__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5379__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8317__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5551__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6659__B _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6500__A1 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8843__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8253__A1 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7950_ _0715_ _1623_ _3304_ _3157_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6901_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7002__C _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7881_ _3196_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8556__A2 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _1376_ _1311_ _2239_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_39_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6763_ _1770_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8308__A2 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8502_ _3789_ _0544_ _2446_ _3791_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5714_ _1239_ _4118_ _1242_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6319__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6694_ as2650.stack\[4\]\[6\] _2134_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5790__A2 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7953__B _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8433_ _3735_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8364_ _3028_ _3567_ _2664_ _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5576_ _1115_ _1121_ _1124_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7315_ _2678_ _2360_ _2688_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4527_ as2650.carry _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7819__A1 _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8295_ _1647_ _0886_ _3603_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7244__I _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7295__A2 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8492__A1 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7246_ _2616_ _2619_ _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4458_ _4038_ _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ as2650.cycle\[5\] _2556_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A4 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4389_ _3969_ _3936_ _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _1548_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7047__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A1 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8075__I _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6059_ _1291_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__A1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4536__C _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8716__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5781__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6089__A3 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8483__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6993__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8235__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7038__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5049__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7210__A2 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5772__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _0963_ _0984_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4688__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4878__A4 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7100_ _1544_ _3950_ _2484_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _3891_ _3892_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8080_ _1322_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8474__A1 _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _0336_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5288__B2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7031_ _4215_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5312__I _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7933_ _1528_ _3287_ _3288_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8739__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7667__C _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7864_ _1632_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _2219_ _1734_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7201__A2 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7795_ _3150_ _4183_ _3151_ _3154_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6960__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4799__S _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4971__B1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6677_ as2650.stack\[4\]\[1\] _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5982__I _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8498__C _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8416_ _2259_ _1297_ _3700_ _2817_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6712__A1 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5515__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ _1170_ _1161_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8347_ _3903_ _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5559_ _3998_ _1101_ _1102_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8465__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8278_ _2407_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5279__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7229_ _2604_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7440__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__A1 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8201__C _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8456__A1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8208__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5442__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5442__B2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4930_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4861_ net8 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6600_ _1974_ _2051_ _2012_ _2013_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5745__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7580_ _2903_ _2909_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4792_ _4073_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6898__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6531_ _1923_ _1925_ _1941_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6462_ _1872_ _1893_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8201_ _3485_ _3512_ _3513_ _3135_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5413_ _0943_ as2650.stack\[5\]\[9\] as2650.stack\[4\]\[9\] _0968_ _0969_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6393_ _1811_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6170__A2 _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8132_ _2734_ _3424_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8447__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5344_ _0896_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6458__B1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8063_ _1614_ _3378_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5275_ _0415_ _0613_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7014_ _2375_ _2282_ _2409_ _3932_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5681__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5433__A1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7916_ _3266_ _0586_ _3272_ _1643_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7186__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7847_ _2471_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6933__A1 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7778_ as2650.pc\[14\] _3139_ _2497_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6729_ _2157_ _0956_ _2160_ _4216_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_109_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7489__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8438__A1 _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6449__B1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7110__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6048__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7413__A2 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5887__I _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4791__I _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A1 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _0618_ _0619_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_42_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__A1 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4466__A2 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6612__B1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8173__I _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8750_ _0149_ clknet_3_5_0_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _1201_ _1465_ _1470_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5966__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7701_ _3009_ _3052_ _2623_ _2495_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _0471_ _0369_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7168__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8681_ _0080_ clknet_leaf_25_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ _1415_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7632_ _2916_ _2996_ _2999_ _2666_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4844_ _0309_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5718__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7563_ _2794_ as2650.stack\[1\]\[6\] as2650.stack\[0\]\[6\] _2789_ _2933_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4775_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6391__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6514_ _1916_ _1945_ _1967_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7494_ _2852_ _2864_ _2767_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _4271_ _1821_ _1850_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7340__A1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6376_ _1832_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4876__I _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8115_ _3428_ _3429_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5327_ _4239_ _0864_ _0867_ _4059_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_114_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8046_ _3326_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5258_ _0782_ _0794_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4457__A2 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _3939_ _0714_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5406__A1 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__S1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8879_ _0278_ clknet_leaf_60_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7427__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A1 _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7331__A1 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7882__A2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4696__A2 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4786__I _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5893__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7162__I _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7634__A2 _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4448__A2 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7398__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8207__B _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__B _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7765__C _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7570__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _4138_ _4139_ _4140_ _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _4071_ _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__A1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__B1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _1164_ _1467_ _1710_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ _4069_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7072__I _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _4103_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7625__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _3991_ _4195_ _1397_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _0506_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7800__I _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7389__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__B _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8802_ _0201_ clknet_leaf_20_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8050__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6994_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5939__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6061__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8733_ _0132_ clknet_leaf_44_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _1449_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8664_ _0063_ clknet_leaf_32_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _1271_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7615_ as2650.pc\[8\] _1536_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _3976_ as2650.idx_ctrl\[0\] _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7561__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8595_ _3242_ _3877_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4375__A1 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7546_ _2500_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4758_ _0318_ _0319_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6116__A2 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7313__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7477_ _1152_ _2607_ _2848_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4689_ _4268_ _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _4254_ _0826_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5875__A1 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _1809_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8029_ as2650.stack\[4\]\[8\] _2134_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8041__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7552__A1 _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7552__B2 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7855__A2 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5866__A1 _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7106__B _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8622__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8032__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__B _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8772__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _1263_ _3961_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5661_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7400_ _1144_ _1138_ _1129_ _2673_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4612_ _3958_ _4155_ _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8380_ _3626_ _3628_ _2216_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5592_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7331_ _2665_ _2663_ _2672_ _2694_ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _4122_ _3905_ _4123_ _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7262_ _1591_ _2361_ _2612_ _1729_ _2637_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__7846__A2 _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4474_ _4054_ _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5857__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ as2650.stack\[0\]\[6\] _1449_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7193_ _2355_ _2570_ _2544_ _2515_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _4142_ _0529_ _1637_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_135_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5609__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8271__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6282__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5085__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ _4079_ _0586_ _4093_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _2368_ _2371_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7782__A1 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8716_ _0115_ clknet_leaf_64_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4596__A1 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ as2650.r123_2\[3\]\[7\] _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8647_ _0046_ clknet_leaf_71_wb_clk_i as2650.r123_2\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5859_ _0438_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4348__A1 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8578_ _2251_ _2433_ _3854_ _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4899__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7529_ _2898_ _2850_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7705__I _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8645__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8795__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8014__A2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7773__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7525__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5839__A1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8253__A2 _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7350__I _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6394__C _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6264__A1 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6900_ _1611_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7880_ _3197_ _3229_ _3237_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_63_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7064__I0 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6831_ _1082_ _1084_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7764__A1 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6567__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__A1 _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6762_ _2113_ _2151_ _2161_ _1060_ _2187_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_108_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8501_ _3790_ _1426_ _3789_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6319__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6693_ _1172_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8432_ _4186_ _4198_ _3734_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5644_ _1183_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8363_ _3028_ _2283_ _3562_ _3669_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5575_ as2650.stack\[5\]\[0\] _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7314_ _4271_ _2633_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4526_ _4106_ _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7819__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8668__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8294_ _3574_ _3578_ _3602_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ _4036_ _4037_ _3994_ _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8492__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _2553_ _2554_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4388_ _3925_ _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8244__A2 _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5058__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _1362_ _1381_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _0411_ as2650.r123\[1\]\[5\] _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7055__I0 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4833__B _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__A1 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6558__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__A1 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5230__A2 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7507__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8180__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8483__A2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7038__A3 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5049__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A1 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7773__C _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__B2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8810__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6182__B1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6721__A2 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__A1 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5360_ _0915_ _0916_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4311_ as2650.ins_reg\[1\] _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5291_ _0844_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8474__A2 _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5288__A2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7030_ _1385_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__A2 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7932_ _1684_ _1361_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7948__C _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _3208_ _3209_ _3218_ _3219_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _1311_ _1084_ _2220_ _2222_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7794_ _1318_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6745_ _2157_ _1018_ _2160_ _1005_ _2166_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6960__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__B2 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _2120_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8415_ _3701_ _3688_ _2261_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5627_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6712__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5515__A3 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8346_ _3388_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4723__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5558_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4509_ _4089_ _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8277_ _3425_ _3586_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8465__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5489_ as2650.stack\[3\]\[13\] as2650.stack\[0\]\[13\] as2650.stack\[1\]\[13\] as2650.stack\[2\]\[13\]
+ _1014_ _1015_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7228_ _2316_ _2317_ _2589_ _2603_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_104_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8086__I _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7159_ _3984_ _2517_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8217__A2 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6228__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7425__B1 _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6779__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7976__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8035__B _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8833__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6951__A2 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8153__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7165__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7900__A1 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6703__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8208__A2 _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5442__A2 as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7195__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7784__B _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _4071_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ _1929_ _1983_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8144__A1 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4699__I _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _1866_ _1896_ _1915_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7075__I _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8200_ net31 _3389_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5412_ _0945_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6392_ _0659_ _4251_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8131_ _3443_ _3445_ _3281_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _0494_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8447__A2 _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7803__I _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8062_ _0851_ _1597_ _1616_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5274_ _0416_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7013_ _2319_ _3972_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5681__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8781__D _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6582__C _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8856__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7915_ _3160_ _3270_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7846_ _3205_ _4244_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8383__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7186__A2 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_77_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7777_ as2650.pc\[13\] _3110_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6394__B1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6933__A2 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ _0543_ _0450_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4944__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6728_ _2153_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8135__A1 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6659_ _1175_ _1853_ _1815_ _2108_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6697__A1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8329_ net35 _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8438__A2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6757__C _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7110__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5121__B2 _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7949__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6924__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6013__B _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8729__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5360__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7637__B1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8879__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4982__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6612__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6612__B2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ as2650.stack\[1\]\[9\] _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7700_ _1000_ _2752_ _3052_ _3065_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_93_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _0464_ _4189_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8680_ _0079_ clknet_leaf_24_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5892_ _0895_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7168__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8365__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7631_ _2630_ _2461_ _2997_ _2998_ _2521_ _2632_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_4843_ _0397_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8403__B _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7562_ _2533_ _2924_ _2931_ _1735_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4926__A1 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _0318_ _0319_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6391__A3 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6513_ _1918_ _1944_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7493_ _2611_ _2851_ _2861_ _2863_ _2504_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _1814_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7340__A2 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6375_ _3994_ _1816_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8114_ _2250_ _4238_ _4241_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_66_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5326_ _4106_ _0591_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5103__A1 _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8045_ _2116_ _3333_ _3368_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5257_ _0795_ _0813_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5053__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6851__A1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4457__A3 _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5654__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5188_ _3939_ _0714_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_116_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4892__I _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7159__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8356__A1 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8878_ _0277_ clknet_leaf_77_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8356__B2 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7829_ _4119_ _3189_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6906__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__A1 _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5893__A2 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7095__A1 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6059__I _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7095__B2 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7398__A2 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8595__A1 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6950__C _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4471__I3 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8223__B _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7570__A2 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7781__C _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4490_ _3966_ _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7322__A2 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4977__I _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A1 as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6397__C _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6160_ _0558_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5111_ as2650.r123\[1\]\[6\] as2650.r123\[0\]\[6\] as2650.r123_2\[1\]\[6\] as2650.r123_2\[0\]\[6\]
+ _3883_ _3889_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _4196_ _1585_ _1375_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__A1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _0503_ _0508_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8801_ _0200_ clknet_leaf_20_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6993_ _1090_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6061__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8732_ _0131_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5944_ _1217_ _1450_ _1457_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7956__C _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8338__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8663_ _0062_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5875_ _1397_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7528__I _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7010__A1 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7614_ _2620_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4826_ _4226_ _0379_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8594_ as2650.psu\[4\] _3874_ _3876_ _3870_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7561__A2 _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4375__A2 _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7545_ _1170_ _2870_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ as2650.holding_reg\[2\] _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7476_ _2709_ _2846_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6116__A3 _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4688_ net6 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8510__A1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _1880_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5324__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6358_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _4106_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6289_ _1112_ _1480_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6824__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8028_ _2120_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4571__B as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7552__A2 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7882__B _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8501__A1 _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__A3 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5315__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5866__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7106__C _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7068__A1 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6815__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4677__I0 as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__I _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4841__A3 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6961__B net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7240__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6252__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__C _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _0308_ _1158_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _4026_ _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5591_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_117_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7330_ _2654_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4542_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7261_ _1117_ _1728_ _2239_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5306__A1 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4473_ _4047_ _4053_ _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4500__I _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6212_ _1164_ _1452_ _1700_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5857__A2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _0754_ _1506_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6074_ _1278_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6282__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7032__B _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8559__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7686__C _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _1267_ _2360_ _2236_ _2372_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8715_ _0114_ clknet_leaf_66_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5927_ _1445_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4596__A2 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7258__I _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8646_ _0045_ clknet_leaf_46_wb_clk_i as2650.r123_2\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5858_ _1370_ _1375_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4348__A2 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _4250_ _0350_ _0361_ _0371_ _4067_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5789_ _1287_ _1303_ _1320_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8577_ _3860_ _3862_ _2492_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7528_ _2853_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7298__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7459_ _2829_ _2830_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4410__I _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__A2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__B2 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__A2 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7222__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7773__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5784__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7525__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5536__A1 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8501__B _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5416__I _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4320__I _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7461__A1 _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6264__A2 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__A1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6016__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7064__I1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _1731_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5775__A1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ as2650.r123_2\[0\]\[7\] _2151_ _2161_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5712_ _1243_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8500_ _1418_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6692_ _2133_ _2131_ _2135_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6319__A3 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7516__A2 _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8431_ _3731_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5643_ _1081_ _1080_ _1110_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5527__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8362_ _2481_ _3665_ _3032_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7313_ _1091_ _2686_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8477__B1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4525_ _4098_ _4102_ _4105_ _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8293_ _1538_ _0726_ _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _2494_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4456_ _3905_ _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ _2553_ _2554_ _2555_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4502__A2 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4387_ _3967_ _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ _1261_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6157__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _1551_ _1552_ _0869_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ _3892_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5996__I _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A2 _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _3913_ _1288_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7507__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8629_ _0028_ clknet_leaf_20_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8180__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6191__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8612__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7691__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7038__A4 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7443__A1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6246__A2 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6067__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7994__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4315__I _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7626__I _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6182__B2 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4310_ as2650.ins_reg\[0\] _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ _0752_ _0762_ _0750_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8474__A3 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7682__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4496__A1 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6237__A2 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7985__A2 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7931_ _3169_ _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7862_ _4267_ _1721_ _3221_ _1335_ _3202_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_51_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _1094_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _3153_ _4131_ _3150_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _1964_ _2164_ _2174_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8635__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4420__A1 _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _1133_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8414_ net40 _3717_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5626_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8345_ _1190_ _3422_ _3646_ _3652_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5557_ _1103_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4723__A2 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4508_ _4086_ _3894_ _4087_ _4088_ _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8276_ _1541_ _3427_ _3579_ _3432_ _3585_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_104_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _1012_ as2650.stack\[7\]\[13\] as2650.stack\[6\]\[13\] _1007_ _0954_ _1040_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__8465__A3 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6476__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _2374_ _2596_ _2600_ _2602_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_78_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4439_ _4019_ _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7158_ _1285_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__A1 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6228__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__B _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6109_ _1243_ _4191_ _4148_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7089_ _3913_ _1370_ _2473_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__A2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A3 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4411__A1 _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7446__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8153__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7900__A2 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4650__B2 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4790_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4402__A1 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4953__A2 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6260__I _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6460_ _1869_ _1895_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6155__A1 _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _0919_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6391_ _1412_ _1071_ _3962_ _1819_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8130_ _3444_ _2670_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5342_ _4120_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6458__A2 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8061_ _2138_ _3327_ _3377_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ _0504_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7012_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7959__C _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__B1 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5969__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7914_ _3213_ _0370_ _1566_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7845_ _2569_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8383__A2 _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6394__A1 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7776_ _3132_ _3009_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6394__B2 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _4129_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6727_ _4036_ _1081_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4944__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _1360_ _1845_ _2106_ _2107_ _1808_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6697__A2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7894__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _1025_ _1127_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _1899_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8328_ net36 _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7646__A1 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__A2 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8259_ _2898_ _3422_ _3561_ _3453_ _3569_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5514__I _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5121__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7869__C _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7949__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8071__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8800__CLK clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A1 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A2 _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A1 _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6688__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7885__A1 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__A2 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7637__A1 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7637__B2 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5112__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6860__A2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7779__C _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8062__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _1466_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _4176_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5891_ _1416_ _4006_ _3997_ _4203_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7630_ _1729_ _2991_ _2678_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _0398_ _0402_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7561_ _1541_ _2829_ _2928_ _2930_ _2628_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4773_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7086__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _1947_ _1966_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6391__A4 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7492_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7876__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6443_ _1769_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6374_ _0495_ _1810_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7628__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ _0870_ _4066_ _0881_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8113_ _4068_ _4061_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_103_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5256_ _0798_ _0800_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8823__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8044_ as2650.stack\[7\]\[0\] _3335_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6300__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ as2650.holding_reg\[6\] _3939_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8053__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__I _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8877_ _0276_ clknet_leaf_74_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7828_ _4123_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6367__A1 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ _1221_ _2659_ _3122_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__I _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6119__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A3 _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5342__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7095__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6075__I _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5030__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7858__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8846__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _4099_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8283__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _4145_ _1576_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5041_ _0510_ _0509_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__A2 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4926__C _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8035__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8800_ _0199_ clknet_3_7_0_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _1735_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8731_ _0130_ clknet_leaf_46_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5943_ as2650.stack\[0\]\[11\] _1454_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8338__A2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8662_ _0061_ clknet_leaf_22_wb_clk_i as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5874_ _1398_ _1399_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7010__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _1177_ _2849_ _2981_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4825_ _0372_ _0376_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5021__A1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8593_ _3875_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7544_ _1169_ _2870_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _4258_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7849__A1 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4687_ _4262_ _4266_ _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7475_ _2581_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8510__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6426_ _0821_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5324__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _4040_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8274__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ _0446_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6288_ _1179_ _1485_ _1752_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5999__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6824__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8027_ _1123_ _1237_ _3358_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _0499_ _0796_ _0797_ _0699_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__A1 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6588__A1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7785__B1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8929_ net46 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8324__B _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8719__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6623__I _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6760__A1 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8869__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8501__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5315__A2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5866__A3 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6815__A2 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5702__I _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__A1 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4677__I1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8017__A1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4318__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A4 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__A1 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _4002_ _4190_ _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5590_ as2650.pc\[2\] _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6751__A1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4541_ _4121_ _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7260_ _2632_ _2634_ _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4472_ _4050_ _3893_ _4051_ _4052_ _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6503__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5306__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6211_ as2650.stack\[0\]\[5\] _1696_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7191_ _2486_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5857__A3 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _4289_ _0296_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _1547_ _1549_ _1550_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4817__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5024_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8559__A2 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6644__S _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _3932_ _3985_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8714_ _0113_ clknet_leaf_66_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5926_ as2650.r123_2\[3\]\[6\] _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6990__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7983__B _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8645_ _0044_ clknet_3_1_0_wb_clk_i as2650.r123_2\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _1376_ _1377_ _1379_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _4032_ _0370_ _4111_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8576_ _3855_ _3861_ _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ _1321_ _1296_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4898__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ as2650.pc\[6\] _2853_ _2850_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4739_ _4283_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7298__A2 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8495__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7458_ _2825_ _2781_ _2827_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_79_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6409_ _1775_ _1803_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7389_ as2650.pc\[2\] _0351_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8247__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8247__B2 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5522__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4808__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7877__C _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5784__A2 _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6981__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8691__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5536__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7133__B _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5432__I _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7461__A2 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7787__C _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8410__A1 _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7213__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6016__A3 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7359__I _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__A1 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ _2095_ _2163_ _2186_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5775__A2 _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6972__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ as2650.cycle\[7\] as2650.cycle\[6\] _3928_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6691_ as2650.stack\[4\]\[5\] _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8430_ _3732_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5642_ _1078_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5527__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8361_ _3541_ _3658_ _3667_ _3296_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5573_ _1113_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5607__I _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7312_ _2684_ _2685_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8477__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4524_ _4103_ _4104_ _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8292_ _2947_ _3600_ _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7243_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4455_ _3969_ _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8229__A1 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7174_ _2553_ _2554_ _2402_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4386_ _3966_ _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _1574_ _1578_ _1584_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _0741_ _0655_ _0417_ _0366_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_58_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5463__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _3889_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7697__C _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8401__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7269__I _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _3950_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5230__A4 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5909_ _1426_ _1434_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6889_ _1281_ _1250_ _2287_ _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_50_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6901__I _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8628_ _0027_ clknet_leaf_34_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7218__B _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8559_ _2280_ _3846_ _3845_ _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4421__I _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8468__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7691__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7179__I _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5206__A1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5206__B2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6954__A1 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__I1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A1 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6182__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8459__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6967__B _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8474__A4 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__A2 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A1 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6258__I _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4740__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7930_ _3159_ _1351_ _3284_ _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7198__A1 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _3913_ _1098_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4506__I _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5748__A2 _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7792_ _3152_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6945__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ as2650.r123_2\[0\]\[2\] _2165_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4420__A2 _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ _2116_ _2119_ _2122_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _3716_ _3703_ _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5625_ as2650.pc\[6\] _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7370__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5337__I _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8344_ _2656_ _3651_ _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5556_ _4155_ _4100_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4507_ as2650.r123\[1\]\[1\] as2650.r123\[0\]\[1\] as2650.r123_2\[1\]\[1\] as2650.r123_2\[0\]\[1\]
+ _3882_ _4081_ _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7122__A1 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8275_ _3433_ _3583_ _3584_ _3396_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5487_ _0919_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8465__A4 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7226_ _1313_ _2405_ _2601_ _2368_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _3957_ _4018_ _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ _1285_ as2650.cycle\[2\] _1096_ _2456_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_119_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4369_ _3944_ _3946_ _3949_ _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_101_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__A2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6108_ _1380_ _4203_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7088_ _0439_ _1546_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _0561_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8316__C _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6936__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4411__A2 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7361__A1 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A2 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4326__I as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4650__A2 _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6927__A1 _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__I _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7352__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6155__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _0914_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6390_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4996__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7104__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8060_ as2650.stack\[7\]\[7\] _3324_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5272_ _0819_ _0823_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7011_ _1304_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5418__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5418__B2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5969__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8602__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6091__A1 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout51_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7913_ _0615_ _0896_ _2156_ _2842_ _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7844_ _3201_ _3204_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6918__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _1234_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7591__A1 _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__S _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6726_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6657_ _0873_ _1903_ _1843_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6146__A2 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _1152_ _1131_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6588_ _0548_ _1950_ _2040_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8327_ _2564_ _3630_ _3634_ _3398_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5539_ _3929_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8258_ _2863_ _2861_ _3565_ _1736_ _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_106_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _3995_ _1099_ _1604_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_15_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8189_ _2762_ _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6082__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6621__A3 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A2 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A1 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7457__I _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7334__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7885__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7192__I _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5705__I _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8625__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__B _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8775__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _0471_ _0447_ _0467_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7795__C _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5890_ _4204_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _4085_ _4049_ _0305_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7573__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7560_ _2734_ _2929_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4772_ _4190_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6511_ as2650.r123_2\[2\]\[2\] _1948_ _1965_ _1862_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7491_ _2344_ _1733_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _1771_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7876__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5615__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_66_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8112_ _3426_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _4250_ _0715_ _4065_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5639__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8043_ _1500_ _2121_ _3367_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5255_ _0798_ _0800_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _4126_ _0744_ _4038_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8053__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4614__A2 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8876_ _0275_ clknet_leaf_42_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7827_ _2523_ _2342_ _1579_ _3962_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7277__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6367__A2 _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7564__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7758_ _2896_ _3121_ _3040_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6709_ as2650.stack\[3\]\[4\] _2143_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7316__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ _2256_ _3054_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A1 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8648__CLK clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8798__CLK clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8044__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6055__A1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__S0 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7896__B _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7187__I _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7555__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5030__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7307__A1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5636__S _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7858__A2 _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8283__A2 _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _0511_ _0509_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6833__A3 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5170__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8035__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _2296_ _2367_ _2335_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8730_ _0129_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5942_ _1208_ _1450_ _1456_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8661_ _0060_ clknet_leaf_24_wb_clk_i as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5873_ as2650.psl\[7\] _4000_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4514__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7612_ _2896_ _2980_ _2847_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7010__A3 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4824_ _4114_ _0386_ _4116_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8592_ _1025_ _2355_ _3774_ _1535_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5021__A2 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7543_ _1169_ _2899_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4755_ _4253_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4375__A4 _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4780__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7474_ _2807_ _2814_ _2844_ _2845_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7849__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4686_ _4055_ _4264_ _4265_ _4266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6425_ _4096_ _0614_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8510__A3 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6356_ _3925_ _4002_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5307_ _0542_ _0583_ _0673_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6287_ as2650.stack\[2\]\[7\] _1482_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8026_ as2650.stack\[5\]\[14\] _1114_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5238_ _0364_ _0498_ _0612_ _0497_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6824__A3 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8026__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7785__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7785__B2 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8928_ net47 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5260__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8859_ _0258_ clknet_leaf_18_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7537__A1 _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6760__A2 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5571__I0 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5866__A4 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6815__A3 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8017__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8813__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6200__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _4120_ _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ as2650.r123\[1\]\[0\] as2650.r123\[0\]\[0\] as2650.r123_2\[1\]\[0\] as2650.r123_2\[0\]\[0\]
+ _3891_ _4045_ _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7700__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6503__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ _1155_ _1694_ _1699_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7190_ _4037_ _2559_ _2568_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5857__A4 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8476__I _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ as2650.psl\[7\] _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _1562_ _1565_ _1567_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__A2 _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4509__I _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8008__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7767__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6724__I _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _1394_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8713_ _0112_ clknet_leaf_66_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5925_ _1444_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7519__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8644_ _0043_ clknet_3_4_0_wb_clk_i as2650.r123_2\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _1074_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8192__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8575_ _1344_ _2437_ _3832_ _3246_ _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5787_ _3907_ _3915_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7526_ _2605_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4738_ _4039_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7457_ _2634_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4669_ _4237_ _4248_ _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A2 _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _1775_ _1803_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7388_ _2759_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8247__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6339_ _0364_ _0788_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7290__I _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8009_ _2136_ _3345_ _3348_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7058__I0 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__A1 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8836__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6981__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7893__C _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4992__A1 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8183__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5536__A3 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7133__C _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7997__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7749__A1 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8410__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5224__A2 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5775__A3 _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6972__A2 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ _1096_ _3955_ _3909_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6690_ _2120_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8174__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _1063_ _1067_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7921__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8360_ _3391_ _3663_ _3666_ _3588_ _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4735__A1 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7311_ _2684_ _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4523_ as2650.r123\[1\]\[7\] as2650.r123\[0\]\[7\] as2650.r123_2\[1\]\[7\] as2650.r123_2\[0\]\[7\]
+ _3999_ _3890_ _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8291_ _2904_ _3590_ _2948_ _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8477__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7242_ _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _3885_ _4034_ _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8709__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _1281_ _2539_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4385_ _3897_ _3962_ _3965_ _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6124_ _1590_ _1596_ _1603_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _0374_ _4246_ _4214_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ as2650.r123_2\[1\]\[5\] _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6660__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5463__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__I _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8401__A2 _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6412__A1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6957_ _2354_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5908_ as2650.psu\[5\] _1428_ _1431_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6888_ _1412_ _1599_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5839_ _1176_ _1330_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8627_ _0026_ clknet_leaf_20_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6715__A2 _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4702__I _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8558_ _3790_ _2434_ _2432_ _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7509_ _2877_ _2830_ _2878_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8489_ _2576_ _2429_ _2430_ _1425_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__I _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7979__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6651__A1 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__A1 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6954__A2 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8156__A1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5390__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8459__A2 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5390__B2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6890__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4740__I1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7860_ _1687_ _2273_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6811_ _1371_ _1731_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7791_ _2216_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6945__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6742_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8147__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ as2650.stack\[4\]\[0\] _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6158__B1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8412_ net39 _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ _1048_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8343_ _1190_ _3647_ _3650_ _3567_ _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ _4005_ _3943_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6877__C _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _4051_ _4087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8274_ _1539_ _3436_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5486_ _1009_ as2650.stack\[5\]\[13\] as2650.stack\[4\]\[13\] _1037_ _1038_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7122__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _1267_ _1287_ _1731_ _2330_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4437_ _4016_ _4017_ _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7156_ _2319_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8681__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4368_ _3948_ _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _1600_ _1601_ _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7087_ _2457_ _1385_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _1530_ _1531_ _1532_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8386__A1 _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7989_ _1497_ _3333_ _3336_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4411__A3 _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7361__A2 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8310__A1 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6359__I _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4607__I _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6927__A2 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6822__I _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8129__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5438__I _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7352__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5340_ _3944_ _3996_ _4144_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7104__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5271_ _0789_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7010_ _2218_ _2222_ _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6863__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5901__I _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6615__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6091__A2 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7912_ _3267_ _1388_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8368__A1 _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7843_ _4216_ _3203_ _1633_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6918__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7828__I _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6732__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7040__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4929__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _4147_ _0541_ _0545_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7774_ _1226_ _3098_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6725_ _1073_ _0912_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7879__B1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6656_ _0878_ _1847_ _2105_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6587_ _1950_ _2038_ _2039_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_121_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8326_ _2247_ _3633_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5538_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8257_ _2898_ _3567_ _2664_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5469_ _1021_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7208_ _1599_ _0896_ _2342_ _0495_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8188_ _2717_ _3473_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7512__B _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7139_ _2272_ _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_55_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4427__I _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8359__A1 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7031__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5593__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7334__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8531__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7473__I _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5896__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5721__I _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8062__A3 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5877__B _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8253__B _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ _0401_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7573__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4771_ _0324_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5584__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5168__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6781__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6510_ _1949_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7490_ _2856_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7325__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6441_ _1866_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5336__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _1770_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8111_ _2486_ _3921_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7089__A1 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5323_ _0355_ _0873_ _0880_ _0440_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8042_ as2650.stack\[4\]\[14\] _2118_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5254_ _0810_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5185_ _4237_ _0726_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8589__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7261__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6064__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8875_ _0274_ clknet_leaf_38_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7826_ _1324_ _3184_ _2343_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6367__A3 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7757_ _3100_ _3108_ _3120_ _2982_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4969_ _4289_ _0296_ _4298_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5078__I _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6708_ _2128_ _2141_ _2145_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7688_ _2630_ _2681_ _3003_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8513__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__A1 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _1995_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5327__B2 _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__A2 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8309_ _3563_ _3613_ _3617_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6827__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5541__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6055__A2 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5489__S1 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7896__C _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7004__A1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__B1 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7555__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A2 _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7307__A2 _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8504__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8520__C _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4620__I _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7491__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6294__A2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8742__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5451__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6046__A2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6990_ _2374_ _2380_ _2386_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ as2650.stack\[0\]\[10\] _1454_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7378__I _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8338__A4 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5872_ as2650.psl\[6\] _3999_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8660_ _0059_ clknet_leaf_35_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7611_ _2944_ _2955_ _2979_ _2845_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4823_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5557__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8591_ _3754_ _2441_ _3869_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7542_ _2852_ _2911_ _2767_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4754_ _4284_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5309__A1 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7473_ _2495_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4780__A2 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4685_ _4134_ _4135_ _4018_ _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5626__I _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__I _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6424_ _4096_ _0403_ _0614_ _0580_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6355_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7841__I _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6809__A1 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ _4106_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_143_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6286_ _1173_ _1485_ _1751_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__A2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5237_ _0364_ _0611_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8025_ _1123_ _1230_ _3357_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5361__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6824__A4 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ net2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7234__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _3899_ _3945_ _3947_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7785__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8927_ net46 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7288__I _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6192__I _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8858_ _0257_ clknet_leaf_16_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5548__A1 as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7809_ _3160_ _1842_ _3168_ _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__B1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8789_ _0188_ clknet_leaf_36_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8615__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5571__I1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4677__I3 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7225__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7776__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6830__I _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8250__C _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ as2650.ins_reg\[0\] as2650.ins_reg\[1\] _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7700__A2 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A1 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7661__I _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6140_ _1632_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7464__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7464__B2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__B1 as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _0576_ _0578_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7216__A1 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8425__C _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5778__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6973_ _1107_ _2369_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8712_ _0111_ clknet_leaf_68_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5924_ as2650.r123_2\[3\]\[5\] _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8638__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__A1 _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8643_ _0042_ clknet_opt_2_1_wb_clk_i as2650.r123_2\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _0906_ _1380_ _0911_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7836__I _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8192__A2 _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _0363_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8574_ _3855_ _3859_ _1841_ _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5786_ _1318_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7057__B _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7525_ _1160_ _2849_ _2895_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8788__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5950__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__I _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7456_ _2825_ _2781_ _2827_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4668_ _4246_ _4247_ _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6896__B _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _1805_ _1863_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7387_ as2650.pc\[3\] net8 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4599_ _4160_ _4163_ _4179_ _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ _0787_ _1793_ _1794_ _0825_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6269_ _1741_ _1726_ _1719_ _1101_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5466__B1 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8008_ as2650.stack\[6\]\[6\] _3338_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7207__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6915__I _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5769__A1 as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__B1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4435__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4992__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8183__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7694__A1 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7481__I _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7997__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7749__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4432__A1 _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _0953_ _1067_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6185__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7921__A2 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _4064_ _1119_ _1076_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__A2 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7310_ net6 _4082_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4522_ _4087_ _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _3483_ _3598_ _3599_ _3135_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7685__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7241_ _2466_ _2329_ _2465_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4453_ _3924_ _3981_ _4013_ _4033_ _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_89_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5904__I _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ as2650.cycle\[4\] _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4384_ _3964_ _3965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5160__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _1272_ _1604_ _1610_ _1618_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7988__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _1527_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5005_ _0561_ _0562_ _4074_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6956_ _1556_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _1427_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6887_ _1284_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6176__A1 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8626_ _0025_ clknet_leaf_20_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5838_ _1349_ _1364_ _1365_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7373__B1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7912__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8557_ _3842_ _3803_ _3843_ _3844_ _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5769_ as2650.cycle\[7\] _3910_ _1282_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7508_ _2877_ _2830_ _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7125__B1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8488_ _1531_ _3756_ _3772_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7439_ _2808_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7979__A2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6100__A1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8803__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4662__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__B2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__I3 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8156__A2 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__I _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__A1 _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__B2 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4784__B _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ _0437_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4405__A1 _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7790_ _2570_ _4062_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _0992_ _1019_ _1000_ _2171_ _2166_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__A2 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8147__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4803__I _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6672_ _2120_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6158__B2 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8411_ _3104_ _3714_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5623_ _1150_ _1164_ _1166_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8342_ _2529_ _2989_ _3648_ _3649_ _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5381__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5554_ _3963_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7658__A1 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4505_ _4085_ _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5485_ _0944_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8273_ _2084_ _0722_ _3582_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7224_ _3988_ _2284_ _2597_ _2599_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ as2650.ins_reg\[4\] as2650.ins_reg\[6\] as2650.ins_reg\[7\] _4017_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6330__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8826__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7155_ _2455_ _3984_ _2493_ _2537_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4367_ _3947_ _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6106_ _1264_ _1395_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8083__A1 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7086_ _2228_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8083__B2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7830__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _0427_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4644__A1 _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8386__A2 _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6397__A1 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7594__B1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7988_ as2650.stack\[7\]\[13\] _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _1713_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6149__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8609_ _0008_ clknet_leaf_62_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7897__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8310__A2 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8523__C _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8129__A2 _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__I _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4623__I _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6560__A1 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7155__B _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5454__I _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5270_ _0824_ _0825_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6312__A1 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6863__A2 _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8065__A1 _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7812__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7911_ _4036_ _3210_ _1389_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6091__A3 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7842_ _3202_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6379__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6918__A3 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7040__A2 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ _1227_ _2659_ _3134_ _3135_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4985_ _4147_ _0527_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4533__I _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6724_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7879__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7879__B2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ _1647_ _1820_ _1811_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5606_ as2650.pc\[4\] _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6586_ _0556_ _1951_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8325_ _3631_ _3632_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _1082_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5364__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8256_ _3566_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5468_ _0493_ _0989_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ _2538_ _2580_ _2583_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4419_ _3892_ _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8187_ _1315_ _3499_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5399_ _0931_ _0938_ _0948_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_59_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7138_ _1312_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7512__C _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7069_ _1281_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A1 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A3 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__I _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_24_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4443__I _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6790__A1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8531__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8295__A1 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7022__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4353__I _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6781__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _0284_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _1869_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5336__A2 _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6371_ _1391_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8110_ _1315_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8286__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5322_ _0876_ _0354_ _4074_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7089__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8041_ _1497_ _2121_ _3366_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _0780_ _0803_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4847__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5184_ _4066_ _0740_ _0742_ _3924_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8589__A2 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__A2 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__A3 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5111__I2 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8874_ _0273_ clknet_leaf_38_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A2 _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7825_ _1104_ _2337_ _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7756_ _1031_ _2752_ _3107_ _3119_ _3114_ _2271_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_40_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__A1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4968_ _0466_ _0468_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5575__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6707_ as2650.stack\[3\]\[3\] _2143_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7687_ _2784_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7574__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4899_ _4116_ _0460_ _4038_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6524__A1 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6638_ _0586_ _1952_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _2006_ _2021_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5094__I _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8277__A1 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8308_ _1543_ _2460_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5027__C _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6827__A2 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8239_ _0657_ _0682_ _3549_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_65_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6854__S _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7252__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6055__A3 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8694__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8201__A1 _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5015__B2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4829__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7491__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6049__B _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6046__A3 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5940_ _1201_ _1450_ _1455_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5871_ _4100_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5179__I _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7610_ _2953_ _2968_ _2978_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4822_ _0377_ _0379_ _0380_ _0381_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__5557__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6754__A1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8590_ _3867_ _3871_ _3873_ _3870_ _2493_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7541_ _2902_ _2901_ _2910_ _2862_ _2527_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4753_ _4281_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7472_ _2813_ _2835_ _2842_ _2800_ _2843_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6506__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5309__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4684_ _4263_ _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _1791_ _1877_ _1878_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8259__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8259__B2 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6354_ _4024_ _4030_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6809__A2 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _0650_ _0583_ _0674_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ as2650.stack\[2\]\[6\] _1482_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8024_ as2650.stack\[5\]\[13\] _1114_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5236_ _0365_ _0504_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5493__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7234__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8926_ net46 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8857_ _0256_ clknet_leaf_16_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7808_ _4029_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5548__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8788_ _0187_ clknet_3_3_0_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__B2 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7739_ as2650.pc\[11\] _2084_ _3046_ _3101_ _3102_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_71_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8498__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5038__B _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__B1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__I _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8422__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5236__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4747__B1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8489__A1 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7161__A1 _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5011__I1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A2 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _4029_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5475__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__B2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _0581_ _3895_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7216__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__I _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _1082_ _1263_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6975__A1 _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5778__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8711_ _0110_ clknet_leaf_68_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5923_ _1443_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__A2 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8642_ _0041_ clknet_3_5_0_wb_clk_i as2650.r123_2\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6727__A1 _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5854_ _3991_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4805_ _0366_ _3894_ _4087_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8573_ _3246_ _2442_ _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5785_ _3956_ _3987_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4541__I _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7524_ _2709_ _2894_ _2847_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4736_ _4290_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5950__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7455_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7152__A1 _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _3954_ _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ as2650.r123_2\[2\]\[0\] _1830_ _1861_ _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7386_ as2650.pc\[3\] _0423_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4598_ _4173_ _4178_ _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6337_ _0824_ _0827_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5372__I _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8101__B1 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6268_ _1543_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__A1 _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8007_ _2133_ _3345_ _3347_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5219_ _0581_ _4221_ _0707_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ as2650.stack\[0\]\[0\] _1460_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8404__A1 _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5769__A2 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__B2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__I _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8732__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4451__I _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7694__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8882__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6378__I _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5457__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__B _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6406__B1 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5885__C _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8174__A3 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6185__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4361__I _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6997__B _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _4100_ _4101_ _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7134__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7240_ _2609_ _2611_ _2615_ _2527_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ _4022_ _4032_ _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7605__C _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _2538_ _2551_ _2552_ _4037_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4383_ _3963_ _3904_ _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6122_ _3952_ _1614_ _1615_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_opt_1_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _1335_ _1548_ _0445_ _0865_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8605__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5004_ _3967_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__B _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6948__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _2300_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7847__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5906_ _4003_ _1417_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6886_ _2278_ _2285_ _2286_ _1438_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8625_ _0024_ clknet_leaf_27_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5837_ net20 _1354_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7373__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7373__B2 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8570__B1 _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8556_ _1414_ _2523_ _2287_ _2231_ _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ as2650.cycle\[6\] _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7507_ net1 _0577_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _4295_ _4297_ _4298_ _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_136_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7125__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8487_ _1063_ _3773_ _3779_ _3624_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7125__B2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5699_ as2650.pc\[14\] _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7438_ _2759_ _2809_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7369_ _1734_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8362__B _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__B _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7116__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__C _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5678__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6057__B _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8778__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4405__A2 _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6740_ _2170_ _1816_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6504__C _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ _2117_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7355__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6158__A2 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8410_ _3696_ _1540_ _3101_ _3680_ _3102_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_108_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5622_ as2650.stack\[5\]\[5\] _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8341_ _2247_ _2460_ _3506_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5553_ _3959_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ as2650.r0\[1\] _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5118__B1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8272_ _3580_ _3554_ _3581_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5484_ _0655_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7223_ _1291_ _2598_ _1613_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4435_ as2650.ins_reg\[5\] _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6330__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7154_ _2459_ _2520_ _2526_ _2536_ _2454_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4366_ as2650.ins_reg\[7\] _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6105_ _4020_ _1579_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7085_ _1413_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _0353_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7830__A2 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5841__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4644__A2 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7594__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6397__A2 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7987_ _3326_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7577__I _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7594__B2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6938_ _1324_ _2312_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _1413_ _1253_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5097__I _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8608_ _0007_ clknet_leaf_62_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7897__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8539_ _0862_ _1514_ _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4580__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__A2 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7337__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5735__I _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6560__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__A1 _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7155__C _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6312__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8065__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6076__A1 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7812__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__A2 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7910_ as2650.psu\[4\] _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6091__A4 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7841_ _3196_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6918__A4 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ _2414_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4984_ _0516_ _0544_ _0489_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _0900_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _0868_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__7879__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _1114_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6585_ _0594_ _1835_ _1837_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5645__I _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8324_ _1300_ _2104_ _4123_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5536_ _4175_ _1083_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8255_ _2992_ _2666_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _0987_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7500__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ as2650.psu\[7\] _2538_ _2582_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4418_ _3883_ _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8186_ _1533_ _3427_ _3493_ _3432_ _3498_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_120_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _0951_ as2650.stack\[7\]\[8\] as2650.stack\[6\]\[8\] _0940_ _0954_ _0955_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_120_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7137_ _2356_ _2315_ _1626_ _2519_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_115_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8056__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4349_ as2650.cycle\[1\] _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5380__I _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ _2453_ _1607_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4617__A2 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6019_ _1513_ _1514_ _4280_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5290__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7567__A1 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A4 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7319__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6790__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_64_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A2 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5896__A4 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8295__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6386__I _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8047__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__I _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8106__I _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6230__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8816__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6781__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7166__B _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5465__I _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__A1 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _1808_ _1812_ _1815_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _0562_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7089__A3 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8286__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8040_ as2650.stack\[4\]\[13\] _2118_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5252_ _0781_ _0802_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4847__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6296__I _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8038__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5183_ _0741_ _4065_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__A3 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5111__I3 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7549__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6245__B _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8873_ _0272_ clknet_leaf_39_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7824_ _3998_ _1555_ _1806_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6221__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7755_ _3053_ _3109_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4967_ _4286_ _4287_ _4294_ _0346_ _0322_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_75_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6706_ _2126_ _2141_ _2144_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7686_ _2863_ _3050_ _3051_ _2902_ _2527_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4898_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _0738_ _1812_ _1952_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5375__I as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7721__A1 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _2017_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8307_ _3541_ _3601_ _3615_ _1524_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5519_ _0926_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8277__A2 _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6499_ _1662_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8238_ _3520_ _3547_ _3521_ _3548_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__6827__A3 _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5324__B _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8029__A2 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8169_ _3480_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7788__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5263__A2 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7960__A1 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7712__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A1 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__A2 _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6451__A1 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4364__I as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6203__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4821_ _0382_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6754__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7951__A1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7540_ _2904_ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4752_ _4225_ _0303_ _0315_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ _2801_ _2807_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4683_ _3942_ _3989_ _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7703__A1 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6506__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _1795_ _1798_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4517__A1 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8259__A2 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _4008_ _1809_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7467__B1 as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6809__A3 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6284_ _1164_ _1485_ _1750_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8023_ _1123_ _1224_ _3356_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5235_ _0790_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5166_ _0382_ _0715_ _0717_ _4239_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5097_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6442__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8856_ _0255_ clknet_leaf_15_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8195__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ _1564_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8787_ _0186_ clknet_leaf_2_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6745__A2 _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5999_ _1229_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7942__B2 _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7738_ _3020_ _3047_ _3081_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ _2733_ _3027_ _3035_ _2467_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4508__A1 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7170__A2 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5181__A1 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5833__I _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__A1 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8661__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__A3 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8422__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5236__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_22_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8186__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8186__B2 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7709__B _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__B _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7933__A1 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4747__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__B2 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8489__A2 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7697__B1 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7161__A2 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5172__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5020_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A1 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__B2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6971_ _2332_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6975__A2 _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8710_ _0109_ clknet_leaf_67_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5922_ as2650.r123_2\[3\]\[4\] _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4986__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8177__A1 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4450__A3 _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8641_ _0040_ clknet_3_5_0_wb_clk_i as2650.r123_2\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5853_ _4174_ _4195_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6727__A2 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4804_ as2650.r123\[1\]\[3\] as2650.r123\[0\]\[3\] as2650.r123_2\[1\]\[3\] as2650.r123_2\[0\]\[3\]
+ _3882_ _4081_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4738__A1 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5784_ _1243_ _4008_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8572_ _3856_ _3858_ _2492_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _2851_ _2865_ _2893_ _2845_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _4292_ _4294_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7454_ _0558_ _0412_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4666_ _4245_ _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7152__A2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _1828_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7385_ _2757_ _2710_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4597_ as2650.holding_reg\[0\] _4174_ _4176_ _4177_ _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6336_ _0497_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8684__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8101__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8101__B2 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6267_ _1740_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5218_ _0697_ _0775_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8006_ as2650.stack\[6\]\[5\] _3342_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _1692_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8404__A2 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _0704_ _0707_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_85_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6415__A1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8168__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8839_ _0238_ clknet_leaf_34_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7915__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7143__A2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7264__B _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5154__A1 _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7711__C _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7603__B1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__A2 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4642__I _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6997__C _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _3889_ _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7134__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7174__B _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4451_ _4031_ _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7170_ _1285_ _1633_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4382_ as2650.ins_reg\[3\] _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _0850_ _1598_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_113_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6052_ _0738_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _0543_ _0563_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8398__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__A2 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A1 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6954_ _2335_ _2339_ _2351_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ net24 _2278_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5648__I _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8624_ _0023_ clknet_leaf_30_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ _1361_ _1329_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7373__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8570__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8570__B2 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8555_ _2279_ _2255_ _1431_ _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7506_ _0559_ _0412_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4718_ _4167_ _4168_ _4152_ _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7125__A2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8322__A1 _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5698_ _0786_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8486_ _3773_ _3778_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7084__B _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7437_ _2715_ _2716_ _2760_ _2763_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4649_ _4228_ _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5383__I _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6884__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _2733_ _2740_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6319_ _0869_ _4222_ _0835_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7299_ _2669_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6636__A1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5439__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_18_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5332__B _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8389__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6942__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7061__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5558__I _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8313__A1 _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7116__A2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8313__B2 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__I _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__C _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6852__I _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__B _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _2118_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7355__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1122_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8340_ _2471_ _3639_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5552_ _4170_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8304__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4503_ _4083_ _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5118__A1 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8271_ _3575_ _0653_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5483_ as2650.r123\[0\]\[5\] _0987_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4434_ _4014_ _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7222_ _1575_ _1592_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7153_ _2528_ _2535_ _1688_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4365_ _3945_ _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6104_ _0851_ _1261_ _1598_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_99_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7084_ _2464_ _2468_ _2392_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _4272_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8722__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7043__A1 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7986_ _1494_ _3333_ _3334_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7594__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _2311_ _2318_ _2327_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_74_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _2267_ _2248_ _2269_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8543__A1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8607_ _0006_ clknet_leaf_58_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5819_ _1325_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ as2650.r123\[3\]\[4\] _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8538_ _0747_ _1518_ _3824_ _3825_ _3826_ _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8469_ _1412_ _1273_ _1733_ _1280_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_124_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6857__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7542__B _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7282__A1 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7034__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4399__A2 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7008__I _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8745__CLK clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4323__A2 _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__I as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8065__A3 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7273__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7273__B2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7025__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7025__B2 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7840_ _3156_ _3200_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6379__A3 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7771_ _2496_ _3130_ _3133_ _3123_ _3011_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6784__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6722_ as2650.r123_2\[0\]\[0\] _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8525__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _2076_ _2098_ _2101_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_137_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5604_ _1115_ _1148_ _1149_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _2030_ _2035_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8323_ _1300_ _2104_ _3605_ _3582_ _3606_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_5535_ as2650.ins_reg\[3\] _3958_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8254_ _2898_ _2297_ _3562_ _3564_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _1005_ _0914_ _1018_ _1019_ _0958_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4417_ _3997_ _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7205_ _2581_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5511__A1 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8185_ _3433_ _3496_ _3497_ _3396_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5397_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4348_ as2650.cycle\[7\] as2650.cycle\[6\] _3928_ _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7136_ _1269_ _2518_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7264__A1 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7067_ _1437_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6018_ _1505_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7016__A1 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7969_ _3203_ _3320_ _3322_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8618__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8516__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5050__I0 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4896__B _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_33_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__I _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5502__A1 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8087__C _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7558__A2 _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5746__I _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4544__A2 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5320_ _0736_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7494__A1 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _0774_ _0805_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6297__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _0667_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8872_ _0271_ clknet_leaf_39_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4480__A1 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7549__A2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7823_ _1271_ _1587_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_64_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6757__B1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6221__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7754_ _2497_ _3117_ _2629_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _0518_ _0521_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6705_ as2650.stack\[3\]\[2\] _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5656__I as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7685_ as2650.pc\[10\] _3014_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4897_ _4129_ _0429_ _0449_ _4128_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6636_ _0733_ _1848_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5732__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _2018_ _1977_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7871__I as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8306_ _3441_ _3614_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5518_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _4260_ _0358_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7092__B _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6288__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8237_ _0560_ _0593_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5449_ _1003_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8168_ _2353_ _3476_ _3481_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7237__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7119_ _2357_ _2498_ _2502_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8099_ _3404_ _3414_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5248__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7788__A2 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7111__I _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5566__I _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7228__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__B1 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7779__A2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__I _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8561__B _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _0337_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7951__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4751_ as2650.r123\[1\]\[1\] _4212_ _0314_ _4217_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5962__A1 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ _4091_ _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7470_ _2837_ _2838_ _2841_ _0972_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__7703__A2 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6421_ _1795_ _1798_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5714__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__A2 _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6352_ _3925_ _1070_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5190__A2 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ _0855_ _0859_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_89_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6283_ as2650.stack\[2\]\[5\] _1746_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8022_ as2650.stack\[5\]\[12\] _3352_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5234_ _0705_ _0791_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_97_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A1 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _0377_ _0719_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5096_ net1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4555__I as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6442__A2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A1 _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8855_ _0254_ clknet_leaf_16_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8195__A2 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7806_ _4222_ _3162_ _3163_ _2652_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_77_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8786_ _0185_ clknet_3_3_0_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5402__B1 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5998_ _1494_ _1495_ _1496_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7737_ _3043_ _3080_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5953__A1 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _0309_ _0406_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5386__I _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ _2501_ _3030_ _3034_ _2666_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6619_ _0654_ _1858_ _2070_ _1910_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7599_ _2529_ _2961_ _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_125_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8806__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8365__C _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7225__A4 _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7630__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8186__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6197__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5944__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7697__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7697__B2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7161__A3 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5711__A4 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7449__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8556__B _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8275__C _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__A1 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _2283_ _1276_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5921_ _1442_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8177__A2 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8640_ _0039_ clknet_leaf_38_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5852_ _4200_ _0892_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7924__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6727__A3 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4738__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8571_ _3855_ _3857_ _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5783_ _1310_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7522_ _2864_ _2884_ _2891_ _2800_ _2892_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4734_ _0294_ _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7688__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7635__B _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7453_ _2824_ _0362_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4665_ _4086_ _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6404_ _1831_ _1860_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8829__CLK clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7384_ as2650.pc\[3\] _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4596_ _3941_ _4075_ _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6335_ _0826_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4910__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A1 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6266_ _1739_ _1727_ _1719_ _3998_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7370__B _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8005_ _2130_ _3345_ _3346_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5217_ _0694_ _0710_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6663__A2 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7860__A1 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6197_ _1635_ _1691_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8185__C _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _0579_ _4219_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7612__A1 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5079_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A3 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8838_ _0237_ clknet_leaf_28_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8769_ _0168_ clknet_leaf_14_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__I _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A2 _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5154__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4901__A2 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7851__A1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6675__I _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6406__A2 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7603__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7603__B2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5090__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5754__I _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5145__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4450_ _4023_ _4024_ _4030_ _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_89_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4381_ _3956_ _3961_ _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_125_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6120_ _4015_ _1605_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6645__A2 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6051_ _1546_ _0873_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _0430_ _0431_ _0447_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4408__A1 as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6948__A3 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _2340_ _2347_ _2349_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__4959__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6884_ _2280_ _2283_ _2284_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8623_ _0022_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5835_ _1362_ _1330_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5908__A1 as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8570__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8554_ _1379_ _1382_ _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5766_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8651__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6581__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7505_ _2634_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4717_ _4293_ _4296_ _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8485_ _3070_ _3775_ _3777_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5697_ _1194_ _1230_ _1232_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7436_ as2650.pc\[4\] _0559_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6333__A1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ _4047_ _4053_ _4083_ _4089_ _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_107_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6884__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ _1954_ _2679_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4579_ _4026_ _4159_ _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6318_ _0815_ _0840_ _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7298_ _1116_ as2650.ins_reg\[2\] _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6495__I _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6636__A2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _0353_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4647__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8389__A2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7061__A2 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4743__I _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8010__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8561__A2 _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__B _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8313__A2 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8077__A1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7722__C _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__A2 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7824__A1 _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4653__I _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8674__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8552__A2 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5620_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6563__A1 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _1093_ _1095_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5484__I _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _4080_ _4082_ _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6315__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5118__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8270_ _3575_ _0653_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5482_ _1034_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7221_ _2236_ _2531_ _1086_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4433_ _3933_ _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8068__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7152_ _3986_ _2529_ _2532_ _2534_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4364_ as2650.ins_reg\[6\] _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7815__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _4015_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7083_ _2428_ _2463_ _2465_ _2467_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7204__I _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _4070_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A2 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8240__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7985_ as2650.stack\[7\]\[12\] _3329_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7079__C _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6936_ _1392_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6867_ _2268_ _2245_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8543__A2 _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8606_ _0005_ clknet_3_4_0_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5818_ _1326_ _1347_ _1348_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5357__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6798_ _2211_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8537_ _0648_ _0759_ _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5749_ _3982_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5394__I _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8468_ _1064_ _3164_ _1555_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_108_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7419_ _0917_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8399_ net39 _3703_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4868__A1 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8059__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7806__A1 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A4 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7806__B2 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7114__I _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8697__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8373__C _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7034__A2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__I _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4399__A3 _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__A2 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5348__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8564__B _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5284__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8222__A1 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7025__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6084__B _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7770_ _3131_ _3132_ _2621_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6784__A1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _2150_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8525__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _2077_ _2081_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5339__A2 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A1 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ as2650.stack\[5\]\[3\] _1135_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6583_ _1834_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8289__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8322_ _2247_ _3629_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6103__I _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _4200_ _4000_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8253_ _3563_ _3546_ _2866_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _0913_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _3903_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4416_ _3996_ _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8184_ _0427_ _3436_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5511__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7135_ _3984_ _2517_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4558__I _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4347_ as2650.cycle\[5\] as2650.cycle\[4\] _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7264__A2 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8461__A1 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ _2423_ _2451_ _2452_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5275__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6017_ as2650.psl\[1\] _1502_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8213__A1 _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A1 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5389__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6775__A1 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7968_ _1059_ _3197_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _1291_ _1598_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7818__B _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7899_ _3256_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8516__A2 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5050__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7109__I _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4468__I _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7255__A2 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8384__B _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6616__C _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7019__I _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8559__B _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5250_ _0777_ _0804_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8862__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5181_ _4111_ _0586_ _0735_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7246__A2 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8871_ _0270_ clknet_leaf_41_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5009__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7822_ _3181_ _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6757__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ _2916_ _3112_ _3113_ _3116_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6542__B _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4965_ _0325_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6704_ _1753_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6509__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ _3044_ _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ _0450_ _0451_ _0390_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _1956_ _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1881_ _1978_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5732__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8469__B _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8305_ _1315_ _3611_ _3613_ _3401_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5517_ _3905_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5672__I _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6497_ _1823_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8236_ _1674_ _0593_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5448_ _0988_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8167_ _1139_ _3421_ _3479_ _2661_ _3480_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5379_ _0922_ _0935_ as2650.psu\[2\] _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7237__A2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8098_ _1571_ _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ _0462_ _2423_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6996__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8198__B1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8735__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5971__A2 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7173__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6920__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8379__B _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4931__B1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5582__I _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8425__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7228__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8425__B2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5239__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__A1 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8561__C _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__I _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5962__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7164__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _4260_ _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7972__I _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ _1874_ _1875_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_70_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5714__A2 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5302_ _4147_ _0845_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6282_ _1155_ _1744_ _1749_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8021_ _3350_ _1217_ _3355_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ _0414_ _0400_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7921__B _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8608__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A2 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8416__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5164_ _0456_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _0581_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8758__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5650__A1 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8854_ _0253_ clknet_3_6_0_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8471__C _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7805_ _4108_ _3164_ _3165_ _0902_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8785_ _0184_ clknet_leaf_6_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5402__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ as2650.stack\[2\]\[12\] _1488_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5402__B2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7736_ _3098_ _3099_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4948_ _0373_ _4222_ _0405_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7155__A1 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7667_ _2918_ _3031_ _3022_ _2676_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _0355_ _0422_ _0435_ _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _2068_ _2069_ _1951_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7598_ _2498_ _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6549_ _1990_ _2002_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8219_ _3530_ _3487_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8407__A1 _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8407__B2 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4746__I _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8218__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7630__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5577__I _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6197__A2 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__I _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7792__I _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7697__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7725__C _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5172__A3 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6201__I _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7449__A2 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8556__C _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6076__C _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__A2 _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8572__B _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__I _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5920_ as2650.r123_2\[3\]\[3\] _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5851_ _4196_ _0901_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7385__A1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4391__I _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _0364_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8570_ _1350_ _2437_ _3832_ _3754_ _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5782_ _1313_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _2801_ _2851_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7916__B _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4733_ _4291_ _0296_ _4171_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7137__A1 _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7452_ _0423_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7688__A2 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ _4242_ _4243_ _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6403_ _4183_ _1833_ _1856_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7383_ _1139_ _2607_ _2756_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6360__A2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4595_ _4175_ _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6334_ _1787_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4371__A1 _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _1541_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8004_ as2650.stack\[6\]\[4\] _3342_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7370__C _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _0694_ _0710_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7860__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _1636_ _1690_ _1621_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4566__I _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5147_ _0402_ _0705_ _0706_ _0610_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4426__A2 _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__A1 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8837_ _0236_ clknet_leaf_28_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7376__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5397__I _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7376__B2 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8768_ _0167_ clknet_leaf_7_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7128__A1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ as2650.addr_buff\[3\] _2679_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8699_ _0098_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7117__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6956__I _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7300__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5090__A2 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7367__A1 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7119__A1 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7027__I _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ _3949_ _3960_ _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6866__I _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__A2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1416_ _1256_ _4292_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input7_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5853__A1 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4386__I _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5001_ _4071_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8398__A3 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4408__A2 _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__A4 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _1613_ _1595_ _1065_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _1270_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6883_ _3995_ _2221_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7358__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5834_ _0741_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8622_ _0021_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5908__A2 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ net3 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8553_ _3840_ _3841_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5945__I _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6581__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7504_ _2397_ _2869_ _2874_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4716_ _4084_ _4090_ _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4592__A1 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8484_ _0973_ _2977_ _3776_ _2302_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5696_ as2650.stack\[6\]\[13\] _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7435_ _1151_ _2806_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _4134_ _4135_ _4226_ _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7530__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__A2 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _2734_ _2738_ _2739_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4578_ _3946_ _4144_ _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _0818_ _0839_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7297_ _2667_ _2662_ _2671_ _2614_ _1414_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6248_ _0892_ _1716_ _1724_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4647__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _0559_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7597__A1 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_3_0_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6644__I0 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8397__I0 _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8010__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6324__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7521__A1 _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__A3 _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8387__B _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6686__I _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A2 _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6088__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6627__A3 _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7824__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5835__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7588__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8819__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8001__A2 _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5765__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7760__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _3955_ _1098_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _4081_ _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _1024_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7512__A1 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _2320_ _2489_ _2593_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4432_ _3926_ _4012_ _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5714__B _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7151_ _2282_ _2519_ _2379_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8068__A2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4363_ as2650.ins_reg\[5\] _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7082_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7815__A2 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A2 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7579__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7043__A3 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8240__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7984_ _3324_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _2328_ _2331_ _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6866_ _1241_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8605_ _0004_ clknet_leaf_61_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5817_ net44 _1333_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6797_ as2650.r123\[3\]\[3\] _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7751__A1 _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4565__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _3927_ _3983_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8536_ _0648_ _0759_ _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8467_ _1596_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7418_ _2788_ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8398_ net38 net50 net36 _3638_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_135_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4868__A2 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _2675_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8059__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5817__A1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4754__I _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__A2 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4703__B _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6190__B _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7742__A1 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7733__C _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8641__CLK clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5036__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__B1 _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _0413_ _0419_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8580__B _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__A2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7981__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6720_ _1389_ _1768_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_75_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _2011_ _2099_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7733__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6582_ _0370_ _1844_ _2034_ _1808_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8321_ _3626_ _3628_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7924__B _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5533_ _4204_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8252_ _2391_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _1011_ _1013_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7203_ net4 _2381_ _1582_ _2579_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4415_ _3945_ _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8183_ _0425_ _0459_ _3495_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5395_ _0936_ _0933_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7134_ _1096_ _2456_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4346_ _3908_ _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7065_ _0856_ _2423_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8461__A2 _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6472__A1 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5275__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ _0750_ _1502_ _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7016__A3 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8213__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5027__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6224__A1 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7967_ _2581_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6918_ _1239_ _2312_ _1598_ _2315_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__7818__C _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7898_ _0433_ _1720_ _3220_ _1345_ _3196_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_51_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__B _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6849_ as2650.addr_buff\[2\] _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8519_ _3761_ _3803_ _3805_ _3808_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_87_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__S _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4710__A1 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8664__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6964__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8452__A2 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__I _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4529__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7744__B _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8140__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__I _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7035__I _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4701__A1 _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _4032_ _0738_ _4022_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8443__A2 _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8870_ _0269_ clknet_leaf_64_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A2 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6206__A1 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _1316_ _1603_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6757__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7752_ _2918_ _3114_ _3115_ _2635_ _2219_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4964_ _0522_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ _2123_ _2141_ _2142_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5439__B _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7683_ _3046_ _3048_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7706__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4895_ _4043_ _0444_ _0455_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6634_ _2084_ _1820_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7654__B _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5193__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6565_ _1973_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5732__A3 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8469__C _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8304_ net35 _3612_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4940__A1 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8687__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5516_ _3934_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_121_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _1824_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8131__A1 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8235_ net51 _3545_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5447_ _0396_ _0990_ _0991_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5496__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8166_ _3387_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5378_ _0923_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4329_ as2650.cycle\[5\] as2650.cycle\[4\] _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7117_ _2500_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8097_ _1119_ _3406_ _3411_ _3412_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8434__A2 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5248__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6445__A1 _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7048_ _2258_ _2436_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6996__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8198__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7945__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7945__B2 _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4759__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8370__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8122__A1 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4931__B2 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6684__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7228__A3 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5239__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6987__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7400__A3 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4680_ _4259_ _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8361__A1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5175__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A3 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6350_ _1806_ _3952_ _1768_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8113__A1 _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5301_ _4027_ _0857_ _0858_ _0626_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6281_ as2650.stack\[2\]\[4\] _1746_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5232_ as2650.r0\[5\] _0304_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8020_ as2650.stack\[5\]\[11\] _3352_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5163_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8416__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6427__A1 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4989__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5013__I _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__A3 _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8853_ _0252_ clknet_leaf_15_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7927__A1 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5948__I _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7804_ _1014_ _1387_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8784_ _0183_ clknet_leaf_7_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _1482_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7735_ _1213_ _1205_ _3014_ _1220_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4947_ _0503_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7666_ _2689_ _3032_ _1415_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8352__A1 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4878_ _0438_ _3898_ _3965_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_123_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ _0682_ _1900_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5166__B2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _2502_ _2962_ _2965_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ as2650.r123_2\[2\]\[3\] _1948_ _2001_ _1862_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8104__A1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _1932_ _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6666__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8218_ net31 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7863__B1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8407__A2 _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8149_ _3459_ _3462_ _3433_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6418__A1 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7091__A1 _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8702__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7091__B2 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7918__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4762__I _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8852__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8591__A1 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8343__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8343__B2 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4904__A1 _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6657__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4507__I1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__A3 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5632__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5768__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5850_ _4009_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ as2650.r0\[3\] _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5781_ _1302_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _2886_ _2887_ _2889_ _2890_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4732_ _4293_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7916__C _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7137__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7451_ _2498_ _2822_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6196__I0 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ _4238_ _4241_ _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7688__A3 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6896__A1 _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _4131_ _1858_ _1832_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4594_ _4159_ _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7382_ _2709_ _2755_ _2582_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6333_ _1788_ _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4371__A2 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6264_ _4164_ _1716_ _1738_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5215_ _0690_ _0772_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8003_ _3338_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5320__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8725__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6195_ _1524_ _1640_ _1642_ _1622_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_83_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _4255_ _0401_ _0613_ _4048_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7073__A1 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ _0576_ _0578_ _0582_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5623__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8875__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8836_ _0235_ clknet_leaf_33_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8573__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8767_ _0166_ clknet_leaf_9_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7718_ _3080_ _3082_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8325__A1 _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8698_ _0097_ clknet_leaf_50_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5139__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _1198_ _3015_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6639__A1 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7561__C _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__A2 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4757__I as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__C _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__A1 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5090__A3 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7367__A2 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8564__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8316__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7119__A2 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5550__A1 _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8748__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7827__B1 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4667__I _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5302__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6882__I _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6951_ _1306_ _2296_ _2348_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5902_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6882_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8555__A1 _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8621_ _0020_ clknet_leaf_49_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5833_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8552_ as2650.carry _3838_ _2402_ _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5764_ _4121_ _1283_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8307__A1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7503_ _2728_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4715_ _4137_ _4141_ _4109_ _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8483_ _1063_ _0967_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5695_ _1186_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7434_ _1144_ _2710_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4646_ as2650.idx_ctrl\[1\] _3977_ _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7365_ _2735_ _2686_ _2737_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4577_ _4109_ _4142_ _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8477__C _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ _0809_ _0842_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7296_ _2668_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6247_ _1531_ _1718_ _1719_ _1722_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4647__A3 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6178_ _1656_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7888__I _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5910__B _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ _0602_ _0623_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8546__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8397__I1 _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8819_ _0218_ clknet_leaf_23_wb_clk_i as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6032__I _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_67_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7521__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7572__B _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5871__I _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6875__A4 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7064__S _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6188__B _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4487__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8482__B1 _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7824__A3 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7037__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7588__A2 _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8537__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6548__B1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7466__C _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _4045_ _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5480_ _0599_ _0990_ _0991_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7512__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8578__B _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ _3994_ _4011_ _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ _2383_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4362_ _3942_ _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8068__A3 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6101_ _4024_ _3952_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7081_ _2220_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7579__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__C _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4637__I0 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7983_ _1492_ _3325_ _3332_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6934_ _4121_ _2291_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7657__B _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _1301_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7200__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8604_ _0003_ clknet_leaf_61_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7376__C _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1344_ _1339_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6796_ _2210_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7751__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8535_ _0539_ _0547_ _3821_ _3823_ _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5747_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4565__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8466_ _2170_ _2584_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8488__B _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ _1210_ _1211_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7417_ _2645_ as2650.stack\[5\]\[3\] as2650.stack\[4\]\[3\] _2789_ _2790_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4629_ _4202_ _4209_ _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8397_ _3688_ _3700_ _3701_ _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7348_ _2619_ _2721_ _2621_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7279_ _1119_ _2623_ _2616_ _2641_ _2652_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_85_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__A3 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8519__A1 _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7990__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6190__C _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7742__A2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4556__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8455__B1 _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5106__I _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6481__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__A1 _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6769__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7430__A1 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6233__A2 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__B2 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ _0526_ _0537_ _0540_ _0344_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8580__C _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__B1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7981__A2 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5776__I _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4680__I _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7196__C _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _1059_ _2050_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7733__A2 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__A4 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5601_ _1005_ _1127_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6581_ _1356_ _1903_ _1952_ _2033_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8320_ _3921_ _3627_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5532_ _1071_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8251_ _2330_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _0977_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6400__I _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7202_ _1176_ _2381_ _1582_ _2578_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4414_ _3901_ _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5444__C _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8182_ _3459_ _3460_ _3494_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5394_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7249__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7133_ _2455_ _3930_ _2493_ _2516_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7940__B _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4345_ _3925_ _3904_ _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _1176_ _2267_ _2436_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4855__I _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__A2 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _1510_ _0760_ _0761_ _0751_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7231__I _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7966_ _3310_ _3319_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _2313_ _1605_ _2314_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7897_ _3246_ _3247_ _3157_ _3254_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6848_ _1954_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4538__A2 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _0513_ _2074_ _2200_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8518_ _1392_ _2381_ _3806_ _3807_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8449_ as2650.r123\[2\]\[4\] _3741_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8809__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4710__A2 _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7660__A1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6980__I _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6215__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7963__A2 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5974__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__B _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__A2 _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7479__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8140__A2 _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__A2 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4675__I _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7651__A1 as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7051__I _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__B _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6206__A2 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7820_ _1289_ _3175_ _3179_ _3180_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7919__C _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7954__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7751_ _2817_ _1268_ _2832_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4963_ _0464_ _0523_ _0470_ _0484_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6702_ as2650.stack\[3\]\[1\] _1765_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7682_ _3020_ _3047_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4894_ _4125_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7935__B _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5717__A1 _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6564_ _2015_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5193__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8303_ net34 net51 _3545_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5515_ _0335_ _0895_ _0899_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _1817_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4940__A2 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8131__A2 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8234_ net32 _3531_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _0993_ _0966_ _1000_ _0982_ _0983_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6142__A1 _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8165_ _1137_ _3406_ _3478_ _3412_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7890__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5377_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ _1270_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4328_ _3908_ _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8096_ _2719_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7642__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6445__A2 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7047_ _1344_ _2437_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8198__A2 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7949_ _1739_ _3247_ _3303_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__A1 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8631__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6040__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__C _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8781__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4695__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7228__A4 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7400__A4 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8361__A2 _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8430__I _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6372__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5175__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7046__I _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8113__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5300_ _0856_ _4107_ _0538_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6124__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ _1148_ _1744_ _1748_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5231_ _0783_ _0787_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7872__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4686__A1 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5162_ _0549_ _0715_ _0717_ _4233_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_111_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5093_ _0549_ _0638_ _0649_ _4128_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_112_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__A1 _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8852_ _0251_ clknet_leaf_14_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7803_ _1386_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8783_ _0182_ clknet_leaf_6_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _1223_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7734_ _1219_ as2650.pc\[11\] _3071_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_40_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _0404_ _0506_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_52_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A1 _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8654__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ _2681_ _1091_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4877_ _4020_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8352__A2 _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6616_ _1036_ _1839_ _2036_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6363__A1 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5166__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _2724_ _2951_ _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6547_ _1899_ _2000_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4913__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8104__A2 _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6115__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6478_ _1887_ _1889_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8496__B _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8217_ _3526_ _3527_ _2808_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6666__A2 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7863__A1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5429_ _4283_ _0302_ _0908_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7863__B2 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8148_ _3460_ _3461_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4529__B _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8079_ _2632_ _3394_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4429__A1 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7091__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7918__A2 _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8591__A2 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6035__I _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4601__A1 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8343__A2 _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6354__A1 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5157__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6106__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7854__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5114__I _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__B2 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8677__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _4080_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5780_ _3971_ _3910_ _1294_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _4296_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7137__A3 _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8334__A2 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _2728_ _2815_ _2821_ _2345_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5148__A2 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6345__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ _4238_ _4241_ _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6196__I1 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6896__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7381_ _2712_ _2722_ _2754_ _2656_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4593_ _3941_ _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8098__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6332_ as2650.r0\[6\] _0400_ _0612_ _0414_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6263_ _1428_ _1718_ _1722_ _1737_ _1715_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8002_ _2128_ _3339_ _3344_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5214_ _0693_ _0711_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6194_ _1544_ _1643_ _1686_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ as2650.r0\[2\] _0611_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5024__I _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A2 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _0630_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5084__A1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4831__A1 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8022__A1 as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8835_ _0234_ clknet_leaf_28_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8573__A2 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8766_ _0165_ clknet_3_3_0_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _1184_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7781__B1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _3044_ _3049_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7395__B _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5908__B _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4929_ _0317_ _0470_ _0488_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8697_ _0096_ clknet_leaf_50_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5694__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8325__A2 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7648_ _1189_ _2990_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5139__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__A1 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7579_ _1168_ _2084_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8089__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8261__A1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5075__B2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4773__I _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6811__A2 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A1 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4822__B2 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5090__A4 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8564__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7119__A3 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__A1 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__C _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7827__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7827__B2 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A2 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A3 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6950_ _2281_ _1276_ _1248_ _2159_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4813__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ _0658_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6881_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8620_ _0019_ clknet_leaf_50_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__A2 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5832_ _0676_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6566__A1 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8551_ _3829_ _3831_ _3839_ _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5763_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__A2 _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7502_ _2870_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4714_ _4084_ _4090_ _4293_ _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5447__C _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8482_ _0992_ _2398_ _3774_ _1725_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5694_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6869__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7433_ _1145_ _2607_ _2805_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4645_ _4035_ _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5019__I _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7364_ _2735_ _2686_ _2737_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_85_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4576_ _4154_ _4156_ _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7279__C1 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _0812_ _0841_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7818__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7295_ _2669_ _4270_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6246_ _3885_ _1716_ _1723_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8842__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6177_ _0874_ _0737_ _0442_ _0352_ _0639_ _0657_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _0602_ _0623_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5057__A1 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6254__B1 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4593__I _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _0416_ _4220_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8546__A2 _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8818_ _0217_ clknet_leaf_23_wb_clk_i as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8749_ _0148_ clknet_leaf_54_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5780__A2 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7809__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7285__A2 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8482__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__B2 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8234__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7037__A2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5048__A1 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8537__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8715__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__A1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5771__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _3995_ _3998_ _4003_ _4010_ _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_144_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6720__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _3899_ _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6100_ _1591_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7080_ _1271_ _2310_ _2321_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8473__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6893__I _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _3961_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8225__A1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6787__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7982_ as2650.stack\[7\]\[11\] _3329_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__B2 as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4637__I1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _1732_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7657__C _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6864_ _0730_ _2248_ _2266_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6539__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8603_ _0002_ clknet_leaf_60_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5815_ _1345_ _1340_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7200__A2 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6795_ as2650.r123\[3\]\[2\] _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7229__I _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5211__A1 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8534_ _3822_ _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5746_ _1069_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5762__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8465_ _0438_ _1410_ _2497_ _2369_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_5677_ _1213_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8161__B1 _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7416_ _0935_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4628_ _3924_ _4013_ _4208_ _4125_ _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8396_ _2259_ _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7347_ _4010_ _2712_ _2718_ _2720_ _2392_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_102_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _4135_ _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8464__A1 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7278_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5278__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6229_ as2650.stack\[1\]\[5\] _1706_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6778__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5450__A1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8519__A2 _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5753__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6950__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6978__I _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5882__I _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4498__I _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8455__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__B2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8207__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4492__A2 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6769__A1 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5122__I _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__B _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7194__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ _1145_ _1131_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6580_ _2031_ _1846_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _0945_ _1066_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5792__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8250_ _3541_ _3544_ _3560_ _3296_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7497__A2 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ as2650.stack\[3\]\[11\] as2650.stack\[0\]\[11\] as2650.stack\[1\]\[11\] as2650.stack\[2\]\[11\]
+ _1014_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_7201_ as2650.psu\[7\] _2267_ _2577_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4413_ _3993_ _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8181_ _1663_ _0389_ _0392_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5393_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7132_ _2496_ _2510_ _2514_ _2515_ _2454_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7249__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4344_ _3890_ _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7063_ _2450_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6014_ _0519_ _0539_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6128__I _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7965_ _0878_ _3198_ _1623_ _1624_ _3318_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5967__I _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6916_ _1103_ _1072_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7896_ _3158_ _1351_ _3253_ _1550_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5983__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _2251_ _2246_ _2254_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _2001_ _2191_ _2195_ as2650.r123_2\[1\]\[3\] _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6932__A1 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8517_ _1841_ _2273_ _1566_ _2301_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5729_ _3963_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7488__A2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8448_ _4217_ _2029_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5499__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8379_ _2630_ _2252_ _1297_ _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8437__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5671__A1 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4781__I _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7297__C _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6923__A1 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6151__A2 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8428__A1 _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5561__B _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7100__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7651__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8600__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__I _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7750_ _3100_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ _0429_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5965__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _1756_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7681_ _1196_ _1537_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7167__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4893_ _4043_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _0728_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7935__C _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5717__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _2010_ _2014_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8302_ _1543_ _3426_ _3604_ _3431_ _3610_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ _0932_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6494_ _1769_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4940__A3 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8233_ _2856_ _3543_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7951__B _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5445_ _0994_ _0996_ _0998_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__8419__A1 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8164_ _2505_ _2718_ _3408_ _3477_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8419__B2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _0932_ _0925_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7890__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7115_ _2310_ _2321_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4327_ as2650.cycle\[3\] as2650.cycle\[2\] _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8095_ _2505_ _2612_ _3408_ _3410_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7242__I _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _2376_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5405__A1 _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8073__I _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _1567_ _1624_ _3302_ _1528_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4534__C _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7879_ _1953_ _3198_ _1623_ _4261_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A1 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5708__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6381__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7330__A1 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4695__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5892__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5381__B _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4447__A2 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7397__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5400__I _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4383__A1 _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7321__A1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__B2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ _0497_ _4048_ _0788_ _0785_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4686__A2 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _4226_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _0390_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__A2 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8851_ _0250_ clknet_leaf_15_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7802_ _0912_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8782_ _0181_ clknet_leaf_3_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ _1492_ _1483_ _1493_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7733_ _1213_ _2659_ _3097_ _2415_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _0366_ _4219_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__A2 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4876_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7664_ _1197_ _3015_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8352__A3 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _1844_ _2065_ _2066_ _1995_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7595_ _2378_ _2944_ _2963_ _2344_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7560__A1 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6546_ _0492_ _1833_ _1999_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6477_ _1797_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5980__I _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8216_ _3526_ _2808_ _3527_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5428_ _0965_ _0966_ _0981_ _0982_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5913__C _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ as2650.psu\[1\] _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8147_ _0353_ _0393_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7615__A2 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8078_ _3978_ _4131_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4429__A2 _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6823__B1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7029_ _2420_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7379__A1 _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8040__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7856__B _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4601__A2 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__I _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6354__A2 _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6986__I _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5890__I _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4507__I3 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6935__B _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5093__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__S0 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A1 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ _0286_ _0287_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _4055_ _4239_ _4240_ _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7542__A1 _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6400_ _1824_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4356__A1 as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7380_ _2721_ _2744_ _2751_ _2752_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4592_ _4164_ _4169_ _4172_ _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6331_ as2650.r0\[6\] as2650.r0\[4\] _0399_ _0611_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _4164_ _1736_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5856__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5213_ _0693_ _0711_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8001_ as2650.stack\[6\]\[3\] _3342_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7006__B _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6193_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5144_ _4255_ _0505_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5608__A1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8763__D _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5075_ _0516_ _0544_ _0527_ _0524_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8270__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8621__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__A2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__I _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8834_ _0233_ clknet_leaf_23_wb_clk_i as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8022__A2 _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8765_ _0164_ clknet_leaf_9_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7781__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5977_ _1479_ _1182_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7781__B2 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7716_ as2650.pc\[10\] _2083_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _0489_ _0465_ _4284_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8696_ _0095_ clknet_leaf_25_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _1196_ as2650.pc\[8\] _2990_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7533__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7578_ as2650.pc\[7\] _0727_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8089__A2 _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6529_ _1940_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7297__B1 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5075__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6272__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8013__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__B _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4889__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7827__A2 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8644__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6263__A1 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8794__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8004__A2 _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _1036_ _1385_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6880_ _1415_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8555__A3 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5831_ _1349_ _1358_ _1359_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7763__A1 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7763__B2 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4577__A1 _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5762_ _3907_ _1295_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8550_ _3836_ _3838_ _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7501_ _1160_ _2871_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_6_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4713_ as2650.holding_reg\[1\] _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7515__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8481_ _2354_ _1432_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5693_ _0574_ _1211_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7432_ _2709_ _2804_ _2582_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _4035_ _4185_ _4213_ _4224_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7363_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4575_ _4155_ _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7279__C2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6314_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7294_ _1128_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7818__A2 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5829__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6245_ _1717_ _1718_ _1719_ _1722_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _4201_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8346__I _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5127_ _0316_ _0648_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4874__I _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5057__A2 _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__A1 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__B2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _4085_ _0505_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8817_ _0216_ clknet_leaf_20_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7754__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8081__I _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8748_ _0147_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8679_ _0078_ clknet_leaf_30_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6309__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5780__A3 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8667__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7809__A2 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__A2 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8256__I _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5048__A2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7745__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6548__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__B _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5220__A2 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8170__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__B1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6720__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7335__I _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _3940_ _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8473__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6030_ _1517_ _1523_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8166__I _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8225__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7070__I _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7981_ _1490_ _3325_ _3331_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6787__A2 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4798__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6932_ _4006_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6863_ _2265_ _2245_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8602_ _0001_ clknet_leaf_65_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ _0523_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6794_ _2209_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5211__A2 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8533_ _3815_ _0491_ _0539_ _0547_ _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5745_ _3951_ _1269_ _1277_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8464_ _2992_ _1384_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8161__A1 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5676_ _1125_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8161__B2 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7415_ _2642_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4627_ _3953_ _4021_ _4031_ _4207_ _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_135_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8395_ _3683_ _3684_ _3699_ _3686_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_117_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6711__A2 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7346_ _2719_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _4134_ _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7277_ _2598_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4489_ _4069_ _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5278__A2 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6475__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6228_ _1155_ _1704_ _1709_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8216__A2 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ as2650.psu\[7\] _1299_ _1652_ as2650.psu\[5\] _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_100_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6778__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7975__A1 as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__A1 _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7727__B2 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6950__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6702__A2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6994__I _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput40 net40 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__8455__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4728__B _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6218__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__A3 _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6943__B _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7966__A1 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5559__B _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7194__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8832__CLK clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7493__C _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4952__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ _1063_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4689__I _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5461_ _0916_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7497__A3 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _3988_ _3990_ _3992_ _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7200_ _1301_ _2576_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4704__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5392_ as2650.psu\[2\] _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8180_ _0426_ _0454_ _3492_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_126_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7131_ _1298_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4343_ _3898_ _3923_ _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7249__A3 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8446__A2 _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7062_ _2449_ _0753_ _2421_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ as2650.psl\[1\] _1502_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6209__A1 as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7964_ _1741_ _1643_ _3317_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6915_ _1371_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7709__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7895_ _3213_ _4261_ _3252_ _3169_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6846_ _2252_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8382__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _2198_ _2199_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6932__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8516_ _1720_ _2299_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ _1254_ _1252_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8134__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8447_ _0493_ _3733_ _3745_ _3746_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5659_ _1198_ _1161_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8378_ _3631_ _3632_ _1321_ _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_102_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8437__A2 _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7329_ _2697_ _2699_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6448__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6999__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8705__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5120__A1 _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5671__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7859__B _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7948__A1 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5379__B as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__I _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8373__A1 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4934__A1 _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8125__A1 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4302__I _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8428__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5561__C _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_20_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7100__A2 _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7939__A1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4961_ _0519_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6700_ _2116_ _1763_ _2140_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7680_ _3019_ _2988_ _3045_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7167__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8364__A1 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4892_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6631_ _2076_ _2077_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_60_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4925__A1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6562_ _2010_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4925__B2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8116__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8301_ _3436_ _3608_ _3609_ _3396_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5513_ _1058_ _1062_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6493_ _1829_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4940__A4 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6678__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8232_ _2906_ _3542_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5444_ _0951_ as2650.stack\[7\]\[10\] as2650.stack\[6\]\[10\] _0967_ _0973_ _0999_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8728__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8163_ _2876_ _3472_ _2725_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5350__A1 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ as2650.psu\[2\] _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7890__A3 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7114_ _2497_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4326_ as2650.cycle\[7\] _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8094_ _3400_ _2829_ _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5102__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7045_ _2345_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7947_ _3169_ _3301_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8355__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7878_ _1725_ _1529_ _3157_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6829_ _4279_ _1309_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A2 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6381__A3 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7330__A2 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__A2 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4792__I _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7397__A2 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8594__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8594__B2 _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A2 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8213__B _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7608__I _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4383__A2 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7771__C _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7857__B1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6124__A3 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__B1 _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _0674_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5091_ _0650_ _0583_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8850_ _0249_ clknet_leaf_15_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7801_ _3161_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8781_ _0180_ clknet_3_3_0_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5399__B2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5993_ as2650.stack\[2\]\[11\] _1488_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7732_ _2496_ _3095_ _3096_ _3011_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _4050_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8337__A1 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7663_ _3028_ _3029_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6899__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _0544_ _1845_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7594_ _0876_ _2390_ _2521_ _1241_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6363__A3 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6545_ _0460_ _1858_ _1998_ _1832_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ as2650.r0\[3\] _0826_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8215_ _2760_ _3502_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4877__I _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _0958_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7253__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5874__A2 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8146_ _0389_ _0392_ _1663_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ as2650.psu\[0\] _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4309_ _3889_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8077_ _1530_ _3392_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5289_ _0845_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6823__B2 _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8084__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7379__A2 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8576__A1 _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7428__I _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7551__A2 _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6354__A3 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5562__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4787__I _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6511__B1 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6814__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5411__I _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__A1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5476__S1 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7790__A2 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__I _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _3918_ _4056_ _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4356__A2 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _4171_ _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6330_ as2650.r0\[7\] _0304_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8169__I _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__I _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5305__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _1735_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _2126_ _3339_ _3343_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ _0723_ _0745_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5856__A2 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1256_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5143_ _0698_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_111_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _0630_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6281__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8558__A1 _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8833_ _0232_ clknet_leaf_24_wb_clk_i as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8764_ _0163_ clknet_leaf_1_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _1068_ _1077_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7781__A2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7715_ _1212_ _0728_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4927_ _4292_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8695_ _0094_ clknet_leaf_25_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6152__I _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7646_ _2453_ _3013_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4858_ _0413_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7533__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7577_ _2945_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6741__B1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4789_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6528_ _1979_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A1 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__B2 _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6459_ _1898_ _1914_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A2 _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8129_ _1116_ _4068_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6272__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8549__A1 _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7221__A1 _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A2 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A1 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__A3 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4310__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5838__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7460__A1 _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6263__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ net19 _1354_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5774__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5761_ _3911_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4577__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7500_ _2857_ _2773_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _4291_ _4172_ _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8480_ _1725_ _3756_ _3772_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5692_ _1227_ _1214_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7431_ _2758_ _2768_ _2803_ _2656_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4643_ _4216_ _4217_ _4223_ _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5526__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _0351_ _4252_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4574_ _3996_ _3948_ _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7279__A1 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7017__B _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6313_ _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7279__B2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7293_ as2650.pc\[0\] net5 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5316__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6244_ _1721_ _1310_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _3969_ _1660_ _1665_ _1669_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5126_ _4282_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7451__A1 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5057__A3 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__A2 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ _4256_ _4086_ _0306_ _0403_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5051__I _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__I _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7203__A1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8816_ _0215_ clknet_leaf_33_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8747_ _0146_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4568__A2 _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5959_ _1193_ _1465_ _1468_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8678_ _0077_ clknet_leaf_31_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7506__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7629_ _2313_ _2989_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5517__A1 _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8311__B _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6610__I _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__A1 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5226__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7690__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7442__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__A2 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5756__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4305__I as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8170__A2 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8611__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6181__B2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7681__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8761__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4495__A1 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6395__C _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6236__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7433__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7980_ as2650.stack\[7\]\[10\] _3329_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5444__B1 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6931_ _4008_ _1408_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_48_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _3918_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8601_ _0000_ clknet_leaf_59_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ _0410_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6793_ as2650.r123\[3\]\[1\] _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8532_ _3816_ _3819_ _3820_ _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _1239_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8463_ _3174_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8131__B _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5675_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7526__I _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7414_ _2239_ _2776_ _2786_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4626_ _3970_ _4206_ _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8394_ _3683_ _3075_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7345_ _1413_ _1556_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4557_ _4136_ _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4722__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7276_ _2647_ _2649_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4488_ _4068_ _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6227_ as2650.stack\[1\]\[4\] _1706_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _0935_ _4270_ _0352_ _0932_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8216__A3 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6227__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _0411_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6089_ _1380_ _4195_ _0575_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7975__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__A2 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8634__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_2_1_wb_clk_i clknet_opt_2_0_wb_clk_i clknet_opt_2_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6163__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7372__S _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput30 net30 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7663__A1 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6218__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__C _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7274__S0 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4952__A2 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7346__I _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _0928_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6154__A1 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _3936_ _3991_ _3978_ _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4704__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _0940_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7130_ _2489_ _2513_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _3906_ _3922_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A2 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7061_ _0730_ _2436_ _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7081__I _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _0857_ _1505_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7014__C _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
.ends

