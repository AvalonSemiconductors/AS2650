// This is the unpowered netlist.
module wrapped_as2650 (WEb_raw,
    boot_rom_en,
    bus_cyc,
    bus_we_gpios,
    bus_we_serial_ports,
    bus_we_sid,
    bus_we_timers,
    le_hi_act,
    le_lo_act,
    reset_out,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    RAM_end_addr,
    RAM_start_addr,
    bus_addr,
    bus_data_out,
    bus_in_gpios,
    bus_in_serial_ports,
    bus_in_sid,
    bus_in_timers,
    cs_port,
    io_in,
    io_oeb,
    io_out,
    irq,
    irqs,
    la_data_out,
    rom_bus_in,
    rom_bus_out,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output WEb_raw;
 output boot_rom_en;
 output bus_cyc;
 output bus_we_gpios;
 output bus_we_serial_ports;
 output bus_we_sid;
 output bus_we_timers;
 output le_hi_act;
 output le_lo_act;
 output reset_out;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 output [15:0] RAM_end_addr;
 output [15:0] RAM_start_addr;
 output [5:0] bus_addr;
 output [7:0] bus_data_out;
 input [7:0] bus_in_gpios;
 input [7:0] bus_in_serial_ports;
 input [7:0] bus_in_sid;
 input [7:0] bus_in_timers;
 output [2:0] cs_port;
 input [18:0] io_in;
 output [18:0] io_oeb;
 output [18:0] io_out;
 output [2:0] irq;
 input [6:0] irqs;
 output [55:0] la_data_out;
 input [7:0] rom_bus_in;
 output [7:0] rom_bus_out;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net286;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net265;
 wire net266;
 wire net287;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire \as2650.PC[0] ;
 wire \as2650.PC[10] ;
 wire \as2650.PC[11] ;
 wire \as2650.PC[12] ;
 wire \as2650.PC[1] ;
 wire \as2650.PC[2] ;
 wire \as2650.PC[3] ;
 wire \as2650.PC[4] ;
 wire \as2650.PC[5] ;
 wire \as2650.PC[6] ;
 wire \as2650.PC[7] ;
 wire \as2650.PC[8] ;
 wire \as2650.PC[9] ;
 wire \as2650.chirp_ptr[0] ;
 wire \as2650.chirp_ptr[1] ;
 wire \as2650.chirp_ptr[2] ;
 wire \as2650.chirpchar[0] ;
 wire \as2650.chirpchar[1] ;
 wire \as2650.chirpchar[2] ;
 wire \as2650.chirpchar[3] ;
 wire \as2650.chirpchar[4] ;
 wire \as2650.chirpchar[5] ;
 wire \as2650.chirpchar[6] ;
 wire \as2650.cpu_hidden_rom_enable ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.debug_psl[0] ;
 wire \as2650.debug_psl[1] ;
 wire \as2650.debug_psl[2] ;
 wire \as2650.debug_psl[3] ;
 wire \as2650.debug_psl[4] ;
 wire \as2650.debug_psl[5] ;
 wire \as2650.debug_psl[6] ;
 wire \as2650.debug_psl[7] ;
 wire \as2650.debug_psu[0] ;
 wire \as2650.debug_psu[1] ;
 wire \as2650.debug_psu[2] ;
 wire \as2650.debug_psu[3] ;
 wire \as2650.debug_psu[4] ;
 wire \as2650.debug_psu[5] ;
 wire \as2650.debug_psu[7] ;
 wire \as2650.ext_io_addr[6] ;
 wire \as2650.ext_io_addr[7] ;
 wire \as2650.extend ;
 wire \as2650.indexed_cyc[0] ;
 wire \as2650.indexed_cyc[1] ;
 wire \as2650.indirect_cyc ;
 wire \as2650.indirect_target[0] ;
 wire \as2650.indirect_target[10] ;
 wire \as2650.indirect_target[11] ;
 wire \as2650.indirect_target[12] ;
 wire \as2650.indirect_target[13] ;
 wire \as2650.indirect_target[14] ;
 wire \as2650.indirect_target[15] ;
 wire \as2650.indirect_target[1] ;
 wire \as2650.indirect_target[2] ;
 wire \as2650.indirect_target[3] ;
 wire \as2650.indirect_target[4] ;
 wire \as2650.indirect_target[5] ;
 wire \as2650.indirect_target[6] ;
 wire \as2650.indirect_target[7] ;
 wire \as2650.indirect_target[8] ;
 wire \as2650.indirect_target[9] ;
 wire \as2650.insin[0] ;
 wire \as2650.insin[1] ;
 wire \as2650.insin[2] ;
 wire \as2650.insin[3] ;
 wire \as2650.insin[4] ;
 wire \as2650.insin[5] ;
 wire \as2650.insin[6] ;
 wire \as2650.insin[7] ;
 wire \as2650.instruction_args_latch[0] ;
 wire \as2650.instruction_args_latch[10] ;
 wire \as2650.instruction_args_latch[11] ;
 wire \as2650.instruction_args_latch[12] ;
 wire \as2650.instruction_args_latch[13] ;
 wire \as2650.instruction_args_latch[14] ;
 wire \as2650.instruction_args_latch[15] ;
 wire \as2650.instruction_args_latch[1] ;
 wire \as2650.instruction_args_latch[2] ;
 wire \as2650.instruction_args_latch[3] ;
 wire \as2650.instruction_args_latch[4] ;
 wire \as2650.instruction_args_latch[5] ;
 wire \as2650.instruction_args_latch[6] ;
 wire \as2650.instruction_args_latch[7] ;
 wire \as2650.instruction_args_latch[8] ;
 wire \as2650.instruction_args_latch[9] ;
 wire \as2650.io_bus_we ;
 wire \as2650.irqs_latch[1] ;
 wire \as2650.irqs_latch[2] ;
 wire \as2650.irqs_latch[3] ;
 wire \as2650.irqs_latch[4] ;
 wire \as2650.irqs_latch[5] ;
 wire \as2650.irqs_latch[6] ;
 wire \as2650.irqs_latch[7] ;
 wire \as2650.ivectors_base[0] ;
 wire \as2650.ivectors_base[10] ;
 wire \as2650.ivectors_base[11] ;
 wire \as2650.ivectors_base[1] ;
 wire \as2650.ivectors_base[2] ;
 wire \as2650.ivectors_base[3] ;
 wire \as2650.ivectors_base[4] ;
 wire \as2650.ivectors_base[5] ;
 wire \as2650.ivectors_base[6] ;
 wire \as2650.ivectors_base[7] ;
 wire \as2650.ivectors_base[8] ;
 wire \as2650.ivectors_base[9] ;
 wire \as2650.last_addr[0] ;
 wire \as2650.last_addr[10] ;
 wire \as2650.last_addr[11] ;
 wire \as2650.last_addr[12] ;
 wire \as2650.last_addr[13] ;
 wire \as2650.last_addr[14] ;
 wire \as2650.last_addr[15] ;
 wire \as2650.last_addr[1] ;
 wire \as2650.last_addr[2] ;
 wire \as2650.last_addr[3] ;
 wire \as2650.last_addr[4] ;
 wire \as2650.last_addr[5] ;
 wire \as2650.last_addr[6] ;
 wire \as2650.last_addr[7] ;
 wire \as2650.last_addr[8] ;
 wire \as2650.last_addr[9] ;
 wire \as2650.page_reg[0] ;
 wire \as2650.page_reg[1] ;
 wire \as2650.page_reg[2] ;
 wire \as2650.regs[0][0] ;
 wire \as2650.regs[0][1] ;
 wire \as2650.regs[0][2] ;
 wire \as2650.regs[0][3] ;
 wire \as2650.regs[0][4] ;
 wire \as2650.regs[0][5] ;
 wire \as2650.regs[0][6] ;
 wire \as2650.regs[0][7] ;
 wire \as2650.regs[1][0] ;
 wire \as2650.regs[1][1] ;
 wire \as2650.regs[1][2] ;
 wire \as2650.regs[1][3] ;
 wire \as2650.regs[1][4] ;
 wire \as2650.regs[1][5] ;
 wire \as2650.regs[1][6] ;
 wire \as2650.regs[1][7] ;
 wire \as2650.regs[2][0] ;
 wire \as2650.regs[2][1] ;
 wire \as2650.regs[2][2] ;
 wire \as2650.regs[2][3] ;
 wire \as2650.regs[2][4] ;
 wire \as2650.regs[2][5] ;
 wire \as2650.regs[2][6] ;
 wire \as2650.regs[2][7] ;
 wire \as2650.regs[3][0] ;
 wire \as2650.regs[3][1] ;
 wire \as2650.regs[3][2] ;
 wire \as2650.regs[3][3] ;
 wire \as2650.regs[3][4] ;
 wire \as2650.regs[3][5] ;
 wire \as2650.regs[3][6] ;
 wire \as2650.regs[3][7] ;
 wire \as2650.regs[4][0] ;
 wire \as2650.regs[4][1] ;
 wire \as2650.regs[4][2] ;
 wire \as2650.regs[4][3] ;
 wire \as2650.regs[4][4] ;
 wire \as2650.regs[4][5] ;
 wire \as2650.regs[4][6] ;
 wire \as2650.regs[4][7] ;
 wire \as2650.regs[5][0] ;
 wire \as2650.regs[5][1] ;
 wire \as2650.regs[5][2] ;
 wire \as2650.regs[5][3] ;
 wire \as2650.regs[5][4] ;
 wire \as2650.regs[5][5] ;
 wire \as2650.regs[5][6] ;
 wire \as2650.regs[5][7] ;
 wire \as2650.regs[6][0] ;
 wire \as2650.regs[6][1] ;
 wire \as2650.regs[6][2] ;
 wire \as2650.regs[6][3] ;
 wire \as2650.regs[6][4] ;
 wire \as2650.regs[6][5] ;
 wire \as2650.regs[6][6] ;
 wire \as2650.regs[6][7] ;
 wire \as2650.regs[7][0] ;
 wire \as2650.regs[7][1] ;
 wire \as2650.regs[7][2] ;
 wire \as2650.regs[7][3] ;
 wire \as2650.regs[7][4] ;
 wire \as2650.regs[7][5] ;
 wire \as2650.regs[7][6] ;
 wire \as2650.regs[7][7] ;
 wire \as2650.relative_cyc ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][15] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][15] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][15] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][15] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][15] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][15] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][15] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][15] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][15] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][15] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][15] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][15] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][15] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][15] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][15] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][15] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire \as2650.trap ;
 wire \as2650.warmup[0] ;
 wire \as2650.warmup[1] ;
 wire \as2650.wb_hidden_rom_enable ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_146_wb_clk_i;
 wire clknet_leaf_147_wb_clk_i;
 wire clknet_leaf_148_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_150_wb_clk_i;
 wire clknet_leaf_151_wb_clk_i;
 wire clknet_leaf_152_wb_clk_i;
 wire clknet_leaf_153_wb_clk_i;
 wire clknet_leaf_154_wb_clk_i;
 wire clknet_leaf_155_wb_clk_i;
 wire clknet_leaf_156_wb_clk_i;
 wire clknet_leaf_157_wb_clk_i;
 wire clknet_leaf_158_wb_clk_i;
 wire clknet_leaf_159_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_160_wb_clk_i;
 wire clknet_leaf_161_wb_clk_i;
 wire clknet_leaf_162_wb_clk_i;
 wire clknet_leaf_163_wb_clk_i;
 wire clknet_leaf_164_wb_clk_i;
 wire clknet_leaf_165_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \wb_counter[0] ;
 wire \wb_counter[10] ;
 wire \wb_counter[11] ;
 wire \wb_counter[12] ;
 wire \wb_counter[13] ;
 wire \wb_counter[14] ;
 wire \wb_counter[15] ;
 wire \wb_counter[16] ;
 wire \wb_counter[17] ;
 wire \wb_counter[18] ;
 wire \wb_counter[19] ;
 wire \wb_counter[1] ;
 wire \wb_counter[20] ;
 wire \wb_counter[21] ;
 wire \wb_counter[22] ;
 wire \wb_counter[23] ;
 wire \wb_counter[24] ;
 wire \wb_counter[25] ;
 wire \wb_counter[26] ;
 wire \wb_counter[27] ;
 wire \wb_counter[28] ;
 wire \wb_counter[29] ;
 wire \wb_counter[2] ;
 wire \wb_counter[30] ;
 wire \wb_counter[31] ;
 wire \wb_counter[3] ;
 wire \wb_counter[4] ;
 wire \wb_counter[5] ;
 wire \wb_counter[6] ;
 wire \wb_counter[7] ;
 wire \wb_counter[8] ;
 wire \wb_counter[9] ;
 wire wb_debug_carry;
 wire wb_debug_cc;
 wire wb_feedback_delay;
 wire wb_io3_test;
 wire wb_reset_override;
 wire wb_reset_override_en;
 wire \web_behavior[0] ;
 wire \web_behavior[1] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__I (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05725__I0 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__I (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05731__I0 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05731__S (.I(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__I (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__I (.I(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__A2 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__I (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__A1 (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__A2 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__I (.I(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__A1 (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__I (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I0 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I1 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__S (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__I0 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__I1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__S (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__I0 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__I1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__S (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__I (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__I (.I(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__A2 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__I (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__I (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__A1 (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A2 (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__I (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__I (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__I (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__I (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__I (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__I (.I(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__A1 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__A2 (.I(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__I (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__I (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__I (.I(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__A2 (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__I (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__I (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A1 (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__I (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__I (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A2 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__A1 (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__I (.I(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A3 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__I (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__I (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__I (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__B (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__A1 (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__B (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__B (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__A2 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__A1 (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__B (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A3 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A3 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__B (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__A3 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__I0 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__I1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__A1 (.I(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__A2 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A1 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A2 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A1 (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__A3 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__A1 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__A2 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__B (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__A1 (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__A2 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__A1 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__A2 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__A2 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__A2 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__A2 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A1 (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A2 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__C (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__A2 (.I(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__A2 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A2 (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__I (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__B (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__C (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__I (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__B (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A1 (.I(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__C (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__I (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A2 (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__C (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__A4 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A3 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__A2 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__B2 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A1 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A2 (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__A1 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__C (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__I (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__B (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A1 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__I1 (.I(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__I (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__I (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A1 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__A1 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__C (.I(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__C (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A1 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__I (.I(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__A1 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__I (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__A1 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__I (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__I (.I(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__I (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__B (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__I (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__I (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A2 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A4 (.I(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A2 (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A3 (.I(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__I (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__I (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__I (.I(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__I (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__C (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__I (.I(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__B (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__I (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__I (.I(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__I (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__I (.I(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A2 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__B1 (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__C (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__B (.I(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__I (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I (.I(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__C (.I(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__A1 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__I (.I(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__B (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__C (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__I (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__I (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A2 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__C (.I(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__I (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A1 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A3 (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A4 (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A1 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__A2 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A1 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A2 (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__I (.I(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A1 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A3 (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A1 (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A1 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A2 (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__I (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A4 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__I (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__B2 (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A2 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__A2 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A1 (.I(\as2650.indirect_target[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A2 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A2 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__I1 (.I(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A1 (.I(\as2650.indirect_target[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A2 (.I(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__B1 (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__B2 (.I(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A2 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A4 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__I (.I(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A2 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A2 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__A1 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__A2 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__I (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A1 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A3 (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__I (.I(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__A1 (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__A2 (.I(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A1 (.I(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A2 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__A1 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A2 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A1 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A2 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A2 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A1 (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A2 (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__C (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A2 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__B2 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A3 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A1 (.I(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A2 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A2 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__C (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__A1 (.I(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__I (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A2 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A3 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A1 (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__B2 (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__A3 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A1 (.I(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__A1 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__B2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__A1 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A1 (.I(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A2 (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__A1 (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__A1 (.I(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__A2 (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__B2 (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A1 (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A2 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A3 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__A2 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__A1 (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__A1 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__B2 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__A3 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__B2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A1 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A2 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A3 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A1 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A2 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A1 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A2 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A3 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A2 (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A2 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A1 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__I (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__A1 (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__I (.I(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A2 (.I(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__I (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A1 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__B (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A1 (.I(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A1 (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A2 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A2 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A2 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__B (.I(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A1 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A1 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A1 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A2 (.I(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A2 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A1 (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__C (.I(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__I0 (.I(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__S (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A1 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A2 (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A1 (.I(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A1 (.I(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A2 (.I(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__I (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A1 (.I(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A2 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A2 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A1 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A2 (.I(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__I (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__I (.I(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__B1 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__B2 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A2 (.I(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A4 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A2 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A2 (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__A2 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__B1 (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__I (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__I (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A2 (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__B2 (.I(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__B (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__A3 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A1 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A2 (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A2 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A2 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__I (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__I (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A2 (.I(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__B1 (.I(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__I (.I(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__B2 (.I(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A1 (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__I (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__I (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A2 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A1 (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A2 (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A2 (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A3 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__B2 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__I (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A1 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A1 (.I(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A2 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__B (.I(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A2 (.I(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A1 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A1 (.I(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__B (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A2 (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__A1 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__B1 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__B2 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A1 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A1 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__I (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__B1 (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__B2 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__I0 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__I1 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A1 (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A2 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A2 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__B (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A2 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A1 (.I(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A2 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A1 (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__A1 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__B (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__I (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__I (.I(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__I (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A2 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A3 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A2 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__B (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A2 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A3 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A1 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A2 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__B (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A2 (.I(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__B (.I(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__B2 (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A2 (.I(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A1 (.I(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__I (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__S (.I(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__A1 (.I(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A1 (.I(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__I1 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__I (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__I (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__I (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__I (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__I (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A1 (.I(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__I (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__I (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__I (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__I (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__I (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__I (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__I (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__I0 (.I(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__I1 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__S (.I(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__I (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__I (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__I (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__I (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__I (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__I (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__I (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A3 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__I (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__I (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__I (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__I (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__I (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__I (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__I (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__I (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A1 (.I(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A2 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A1 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A2 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A1 (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__I (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__I (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__I (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__I (.I(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A2 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__I (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__A1 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__A2 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__I (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A2 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A3 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__I (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A2 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__B (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__B (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A2 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__B (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__I (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__I (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__I (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A2 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__I (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A2 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A3 (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__I (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__I (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__I (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__I (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__A4 (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__A1 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__I (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A1 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A2 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__I (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__I (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__I (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A2 (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A3 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__I (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__A2 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__A3 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__I (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__B (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__I (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__I (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A2 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__A2 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__B1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A2 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__I (.I(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__I (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__I (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A2 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__B1 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__I (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A2 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__I (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__I (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__I (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__I (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__I (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__I (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A2 (.I(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A2 (.I(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A2 (.I(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A2 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A2 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__I0 (.I(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__S (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__I0 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__S (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__I (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__A2 (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A2 (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__A2 (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__I1 (.I(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__S (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__I (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__I1 (.I(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A1 (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A2 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__I (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__I (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A1 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A2 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__I (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A2 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A2 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A2 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A1 (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__I (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A4 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A1 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A3 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A1 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__B (.I(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__A2 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__I (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__B (.I(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__I (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A2 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A1 (.I(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__B (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A2 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__I (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A1 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A2 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__I (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A2 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__B (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__I (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__I (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A2 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__B (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__A1 (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A2 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__I (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A2 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__I0 (.I(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__S (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A2 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__I (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__I (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__I (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A2 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__I0 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__S (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__B (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__A1 (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A2 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__I (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__I (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__I (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A2 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__I (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A1 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A2 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__A1 (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A2 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__I (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__I (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A2 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__I (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A1 (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A2 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A1 (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A2 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A2 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A2 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__I (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A1 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A3 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A1 (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A2 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A2 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__I (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A2 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A3 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__I (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A1 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__B (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A2 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A2 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__I0 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__I1 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__I0 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__I1 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__I0 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__I1 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__I0 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__I1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__I0 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__I1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__I0 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__I1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__I0 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__I1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I0 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__I1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__I1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__I1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I0 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__I1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__I1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__I1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__I (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__I1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__I1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__I1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__I1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__I (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__I1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__I1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__I0 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__I1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I0 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__I1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__I (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__I0 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__I1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__I0 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__I1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__I0 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__I1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__I0 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__I1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__I (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__I0 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__I1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__S (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__I0 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__I1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__S (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__I0 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__I1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__S (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__I0 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__I1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__S (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A1 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A2 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A3 (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__I0 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__I1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__S (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__I0 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__I1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__S (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__I0 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__I1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__S (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A2 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__I (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A2 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A2 (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A2 (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__B (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A2 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A1 (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__I (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A2 (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__B (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__I (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A2 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__I (.I(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A1 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A2 (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A1 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A2 (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__B (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A2 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__I (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__I (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__I (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__A2 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__I (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__A1 (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A2 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__B2 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__A1 (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A2 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07077__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__A1 (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A2 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A1 (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A2 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__I (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__I (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__I (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A1 (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A2 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__A1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A1 (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__I (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__I (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A1 (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__I (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A2 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A2 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__I (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__I (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__I (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A1 (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__I (.I(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__I (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__A2 (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__A1 (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__I (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A2 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A1 (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__I (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A2 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A1 (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A2 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A1 (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A2 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__B (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__I (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__C (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A2 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A2 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A2 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__I (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__I (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A1 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A1 (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A1 (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A1 (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__I (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A1 (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A1 (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__I (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__B (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A1 (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__B (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__I (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__B (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__B (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__B1 (.I(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A1 (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__B (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__B (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__B1 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__I (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__B1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A1 (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__B (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__B1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__C (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A1 (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__B (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__C (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A1 (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__B2 (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__B1 (.I(net418));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__C (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A2 (.I(net411));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A3 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__I (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__I (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A1 (.I(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__I (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__B (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A2 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__B (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A1 (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A1 (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__B (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__I (.I(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A2 (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__B (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A1 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A2 (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A1 (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__I (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__I (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A2 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A2 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A2 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A2 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__C (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__B (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__B (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__I (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__B (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A1 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__I (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__I (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__I (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A1 (.I(net87));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A2 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A1 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A3 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A1 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A2 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A2 (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A3 (.I(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A2 (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__I (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A2 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A1 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A2 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A1 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A2 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__I (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A2 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__B1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A1 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A2 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A1 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__C1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__I (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A2 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__B (.I(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A1 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A2 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__B (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A1 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A2 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__I (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__I (.I(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A1 (.I(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A1 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A1 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A2 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A3 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A4 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__I (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A2 (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A3 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A4 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A1 (.I(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A3 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A1 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__B (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A3 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A2 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__C (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__I (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A2 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A2 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__B1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A1 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A2 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__A2 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__I (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__I (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__I (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__I (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__I (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__I (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A2 (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A1 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__I (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A3 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A1 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A2 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__I (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__I (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__I (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A1 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A2 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__I (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__I (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__I (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A2 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__I (.I(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__I (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A1 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A3 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__I (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__S (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__I (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__I (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__I (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A1 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__A1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__A2 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__I (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__I (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__I (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__I (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A2 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A2 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__I (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__S (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__I (.I(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A1 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__I (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__S (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I0 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I1 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A3 (.I(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A2 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A2 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__I (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__I0 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__S (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__S (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__I (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A1 (.I(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A2 (.I(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__I (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A1 (.I(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__I (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__S (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__I (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__I (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A2 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A1 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__I (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__S (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__I (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A1 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A1 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__I0 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__I1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__S (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__I (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__I (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__I (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__I1 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__S (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__I (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__I (.I(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__I (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__I (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A2 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A2 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__I (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__S (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__I (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A1 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A1 (.I(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__I (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A2 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A1 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__S (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A2 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A1 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__S (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__I (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__I (.I(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A1 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A1 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__B (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A1 (.I(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__S (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__I (.I(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__I (.I(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A1 (.I(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A1 (.I(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A2 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__B (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__I (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__I (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A1 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__I (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A1 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__I (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__I1 (.I(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__I (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A2 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__I (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__I (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A2 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__I (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__I (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__I (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__I (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__B (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A1 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__S (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__S (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__S (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__S (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__S (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__S (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__I0 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__S (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__S (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__S (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__S (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__S (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__S (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__I1 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__S (.I(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__S (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__S (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__I0 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__S (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__S (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__S (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__S (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__S (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__S (.I(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__I (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__I1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__I (.I(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A3 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__S (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__S (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__S (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__S (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__I0 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__I1 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__S (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__S (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__S (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__S (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__I1 (.I(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__I1 (.I(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__I1 (.I(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__I1 (.I(\as2650.stack[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__I (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A4 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__I (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__S (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__I (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__I1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__S (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__I (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__S (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__I1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__S (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__I (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__I (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__S (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__I (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__S (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__S (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__I (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__S (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__I (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__S (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__S (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__S (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__S (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__I (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__I (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__I (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__I (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__I (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__I (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__I (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A4 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__I (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__S (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__I1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__S (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__S (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__I1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__S (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__I (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__S (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__S (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__S (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__S (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__I (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__S (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__S (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__S (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__S (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__I (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__S (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__S (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__S (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__S (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__I (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A1 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__S (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__I (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__S (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__I (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__S (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__S (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__I (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__S (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__I (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__S (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__S (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__I (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__S (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__S (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__S (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__S (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__I0 (.I(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__S (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__I (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__I (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__I (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__I (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__I (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A1 (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A3 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__I (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__S (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__I (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__S (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__I (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__S (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__S (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__I (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__S (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__I (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__S (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__I (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__S (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__I (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__S (.I(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__I (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__I (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__S (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__S (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__I (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__S (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__I (.I(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__S (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__I (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__I (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__S (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__I (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__S (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__I (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__S (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__S (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A3 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__S (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__S (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__S (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__S (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__S (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__S (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__S (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__S (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__S (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__S (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__S (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__I1 (.I(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__S (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__I (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__S (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__S (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__S (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__I1 (.I(\as2650.stack[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__S (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A4 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__S (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__S (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__S (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__S (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__S (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__S (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__S (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__S (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__S (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__S (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__S (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__S (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A2 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A4 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__I (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__S (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__I (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__S (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__S (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__S (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__S (.I(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__I (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__S (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__S (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__S (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__S (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__I (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A4 (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__I (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__S (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__S (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__S (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__S (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__I (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__S (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__S (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__S (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__S (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__I (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__S (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__S (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__S (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__S (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__I (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__S (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__S (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__S (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__S (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A1 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__I (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__S (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__S (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__S (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__S (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__I (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__S (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__S (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__S (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__S (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__I (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__S (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__S (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__S (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__S (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__I (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__I0 (.I(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A3 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__I (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__S (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__S (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__S (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__S (.I(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__I (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__S (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__S (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__S (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__S (.I(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__I (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__S (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__S (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__S (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__S (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__I (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__I0 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__S (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__S (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__I1 (.I(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__S (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__S (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__I (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__I (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__I (.I(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A3 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A1 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A3 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A2 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__I (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A3 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__B (.I(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__I (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A1 (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__I (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A2 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A3 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A2 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A1 (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A2 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__I (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A3 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__I (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A1 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A2 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A3 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A2 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A3 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A1 (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A3 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A2 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A4 (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__I (.I(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A2 (.I(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A3 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A1 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A2 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__I (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__A1 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A2 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A3 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A3 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__I (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__S1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__I (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__I (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__I (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__I (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__I (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A1 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A1 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__B (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A1 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A2 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A2 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A2 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A2 (.I(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__I (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__I (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A2 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__I (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__I (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__I (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__B (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__I (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A2 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__I (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__I (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A3 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__I (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A2 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A3 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A4 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__I (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__I (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__B (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__C (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__I (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__I (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__I (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__B1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__I0 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__I3 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__S1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__I (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A1 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__I (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__I (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A2 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__B (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A2 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A1 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__C (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A1 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__B2 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__I (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A1 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A2 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A3 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__B1 (.I(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__C (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__B (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__B (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A1 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__B (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__I (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__I (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__I (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__A1 (.I(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__B1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__I0 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__I1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__I0 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__I1 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__I0 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__I1 (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__S (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A1 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__C (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__I (.I(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__I (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__I (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__I (.I(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__I (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__B (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A1 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__I (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A1 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A1 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A2 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A2 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A4 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A2 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__I (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__I (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__I (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__I (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__I (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__B1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A2 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__I0 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__I1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I0 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__I1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A1 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__A2 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A1 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A2 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A2 (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__I (.I(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__B (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__B (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A1 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A3 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__I (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__I (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__I (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__I (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__I (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__B1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__I (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__I3 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__I0 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__S (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__C (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A2 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A1 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A2 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__I (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A2 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A2 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__I (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__I0 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__I (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__I (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__I (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__I (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__I (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__B1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A2 (.I(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I0 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I3 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A2 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A2 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A1 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__I (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A1 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__A1 (.I(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__I (.I(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__I (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A2 (.I(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__C (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A1 (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A1 (.I(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A1 (.I(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__I (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__I (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__I (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__I (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__B1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__I0 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__I1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A2 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A2 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B2 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__I (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__B (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A1 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__C (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A1 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A2 (.I(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__I (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__I (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A2 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__I (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__I (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__I (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__B1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__I0 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__I1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A2 (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__I (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__I0 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__I1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__S (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__I0 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__I1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__B2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A1 (.I(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__I (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__I (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A2 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__B (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__I (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__I (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__I (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A1 (.I(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__B1 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A2 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__S (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__I0 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__S (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__S (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__I0 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__S (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__S (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__I1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__S (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__S (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__S (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__S (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__S (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__S (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__S (.I(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__I (.I(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__S (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__S (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__S (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__S (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__B (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A2 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A2 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A2 (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__B (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A1 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__B (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__I (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__I (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__I (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__I (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__I (.I(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__I (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__I (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__I (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__I (.I(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__I (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A2 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A3 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A4 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A2 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A1 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__I (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A3 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__B (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A4 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A2 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A3 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A1 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A3 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__I (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A2 (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__I (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A2 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A3 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__B1 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__B2 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__I (.I(\as2650.indirect_target[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__I (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__B (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A2 (.I(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A3 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__B (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__I (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A3 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__I (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__I (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__B2 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__B1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__B2 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A2 (.I(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__B (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__I (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__B1 (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__I (.I(\as2650.indirect_target[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__I0 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__I1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A3 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A2 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__B2 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__B1 (.I(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__B2 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__I0 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__B1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A3 (.I(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__I (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__I (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__B1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__I (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__B1 (.I(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__I (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__I (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__I (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__I (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__I (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A2 (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A2 (.I(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__B1 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__I (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A2 (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A2 (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__B1 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A1 (.I(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__B1 (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__I (.I(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A2 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A1 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__B1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A1 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__I (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A1 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A2 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__B1 (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__B2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__I (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__I (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__I (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A1 (.I(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__B2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A2 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__B (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__I (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A2 (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__I (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A2 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__I (.I(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__I (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__I (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__B2 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__C2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__I (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__B1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__B2 (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__C2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__I (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__I (.I(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A1 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A2 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A3 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A2 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__B2 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__B (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__B2 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__B2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A1 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__I (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__B2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__I (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__I (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A1 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A2 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__B (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__B2 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__B (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A1 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__B (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__B (.I(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__I (.I(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__I (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A1 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A2 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A2 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__I (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__I (.I(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A2 (.I(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A2 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__A2 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__B1 (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A1 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A1 (.I(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A2 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__B1 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__I (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__I (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__I (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__I (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A1 (.I(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A1 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__B (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__I (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A1 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A3 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A1 (.I(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__B (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__I (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A3 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A2 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__B (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__B (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__I (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A1 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A2 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__B (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__B1 (.I(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__B2 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__I (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__B (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A1 (.I(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A2 (.I(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A1 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__I (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__I (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A1 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A2 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__I (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__I (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__I (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__B2 (.I(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A1 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__I (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A1 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A1 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__I (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A1 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__I (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__I (.I(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__B2 (.I(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A1 (.I(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__I (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A1 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__I (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__I (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A2 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A1 (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A2 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__B (.I(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A1 (.I(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__B (.I(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A1 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__B2 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A1 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__B2 (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__I (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__B2 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A1 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__B2 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__B (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__I (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__I (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A1 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A2 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A1 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A2 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__B (.I(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A2 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A3 (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__B2 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__B (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__C (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A3 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A4 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A1 (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__B (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__A4 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__I (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__I (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__B1 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__B2 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__C (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A2 (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A3 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__B2 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__B1 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__C2 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A1 (.I(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__C (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A2 (.I(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A2 (.I(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A1 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A3 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A3 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A1 (.I(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A3 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A4 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__I (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A3 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__I (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__B (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__C (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__B (.I(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__I (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__I (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__I (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__I (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__I (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__I (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__C (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__I (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__C (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A1 (.I(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__I (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__I (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__I (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__I (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__I (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__I (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__I (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__I (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__I (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__C (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__I (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__C (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A2 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__I (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A1 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A2 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__I (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__I (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A2 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A2 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__I (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__I (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__I (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__I (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__I (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__I (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A1 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__B2 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__B2 (.I(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__I (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__I (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__I (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__I (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__B1 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__I (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__I (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__B2 (.I(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__C (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A2 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__B (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__B (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__B (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__C (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A3 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__B (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A3 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A2 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A1 (.I(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A3 (.I(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A1 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A3 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A3 (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A1 (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__B (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A1 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A3 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__I (.I(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A4 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__C (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__C (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A1 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__I (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__I (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__I (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__B1 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__B2 (.I(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A2 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__B1 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__B1 (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__B1 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__B1 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__B2 (.I(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__A1 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__B (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__C (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__C (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__A2 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__I1 (.I(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__I (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__I (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__I (.I(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__B1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__B2 (.I(\as2650.stack[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__B2 (.I(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__B2 (.I(\as2650.stack[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__B1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__B1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__B1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__B1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__B (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__C (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__I (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__I (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__B (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__I (.I(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A2 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__A2 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__B (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A1 (.I(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__I (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A1 (.I(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A1 (.I(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__I (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A1 (.I(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A1 (.I(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A1 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A1 (.I(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__I (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__I (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__I (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__I (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__I (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__B (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A2 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__I (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__I (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__I (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__I (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__I (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__I (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__I (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__I (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__B1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__I (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__I (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__B1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__I (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__I (.I(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__I (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A2 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A1 (.I(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A2 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__S (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__I (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A1 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__I (.I(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__I (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A1 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A1 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__I (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__C (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A1 (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A2 (.I(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__I (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A2 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__B (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__I (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__I (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A2 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A3 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A2 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__A2 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A2 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__I (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__I (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__I (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__I (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__I (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__B1 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__A1 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__I (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A1 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__C (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A1 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__A1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__C (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A3 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__B (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__I (.I(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__I (.I(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__I (.I(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A2 (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__B1 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__I (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__B1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__B1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A2 (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__B1 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__A1 (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A2 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__B1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__B1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__A2 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__B1 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A2 (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__B1 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A1 (.I(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__A2 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A1 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__I (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__B (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__A1 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__C (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__I (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__I (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A1 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A2 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__I (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__B1 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A1 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__I (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A2 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__A1 (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A1 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A2 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__C (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__B (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A2 (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A1 (.I(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A1 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__C (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__C (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A1 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__I (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__I (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__I (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__I (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__I (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__I (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__I (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__I (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A2 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__A1 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__I (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A1 (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__A1 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A1 (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A1 (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__C (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__I (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A3 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__B (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A2 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A1 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__A1 (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A1 (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__A1 (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A2 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A2 (.I(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A1 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A2 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A1 (.I(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__B (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A2 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A1 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__I (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__C (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__I (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__B2 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A1 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A2 (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__B1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__B2 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A2 (.I(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A1 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__B1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__I (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A2 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__A2 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__C (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A1 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A1 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A1 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A2 (.I(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__C (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__B (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__B2 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__C (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__C (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__I (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__I (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A2 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__B1 (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__I (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__I (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__B1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__I (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A2 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__B1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__A2 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__B1 (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__I (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__I (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__B1 (.I(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__B2 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__I (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__I (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A1 (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A2 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__B1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A2 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__B1 (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A1 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__C (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A1 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A2 (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__B (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__I (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A2 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__B (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__A1 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__C (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__C (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__C (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__A2 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__A2 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A2 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__I (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__I (.I(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__I (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A1 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__I (.I(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A1 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A1 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__C (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__I (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__I (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A1 (.I(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A2 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A2 (.I(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A2 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A2 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A2 (.I(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__B1 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__B1 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A2 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__B1 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A2 (.I(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__B1 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A1 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__A1 (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__B (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__A1 (.I(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A1 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A1 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__C (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__C (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A1 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__B (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__C (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A2 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__B1 (.I(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A2 (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__B1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A1 (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__B1 (.I(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__B1 (.I(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A1 (.I(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__B1 (.I(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A1 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A2 (.I(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A3 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A2 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__B (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__C (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A1 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A1 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__A2 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__B (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__B (.I(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__C (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A1 (.I(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__B (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__I (.I(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__A1 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__B1 (.I(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__B2 (.I(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A1 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A3 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__B2 (.I(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__A1 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A1 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A1 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A2 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A1 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__B (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__B (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A2 (.I(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__A1 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__B2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__B (.I(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__B (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__B (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__C (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__I (.I(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__I (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__B1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__I (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__I (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__B1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__B2 (.I(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__B1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__B1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__B1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__B1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__B1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__B1 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__A2 (.I(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A2 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__B (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A1 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__A1 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__I0 (.I(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__A1 (.I(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__B2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__C (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__B (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A1 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__A1 (.I(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__B (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A1 (.I(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__B (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__I (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__I (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__I (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A4 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A2 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A1 (.I(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__A2 (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A2 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__A1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__A2 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A2 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A1 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A2 (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A3 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__A1 (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__A2 (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__I (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__B (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A2 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__B1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__I (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__B (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A1 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__A2 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A2 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A3 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A2 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__I (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__I (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__I (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__I (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A2 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__B (.I(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A2 (.I(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__I (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A2 (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A1 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__I (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__A1 (.I(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__A1 (.I(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__B2 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A1 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__B2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A1 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A1 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__C (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A1 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__A1 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A2 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__A1 (.I(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__B (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A1 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A2 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__B2 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__B2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__I (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__A2 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__B2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__B (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A2 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A2 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__B (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A1 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A2 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A2 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A1 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__A2 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A2 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__A1 (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__A2 (.I(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A1 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A3 (.I(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A3 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A4 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A3 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__B (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__I (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A1 (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__B (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A1 (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__B (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__B (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__B (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__A1 (.I(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__B (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__A2 (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A1 (.I(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A2 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A1 (.I(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__A1 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__B (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A1 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A3 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__I (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A1 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A1 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A2 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A3 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A4 (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A2 (.I(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A4 (.I(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A1 (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__A2 (.I(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__A3 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__A1 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__A3 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__A1 (.I(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__A3 (.I(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A1 (.I(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A3 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__I1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__A1 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A2 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A1 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A3 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A1 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A3 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__A4 (.I(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A2 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A2 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A2 (.I(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A2 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A2 (.I(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A1 (.I(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A2 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__B2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A1 (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A2 (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__B1 (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__A1 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A2 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A1 (.I(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__A1 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__B1 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__B2 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__C1 (.I(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A2 (.I(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__B1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A1 (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A2 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__B2 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A2 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A3 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A4 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A1 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A1 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__A1 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A2 (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__B2 (.I(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__B3 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A1 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A1 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A2 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A1 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A3 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A4 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__I (.I(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A2 (.I(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__A2 (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__A1 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__A2 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__A3 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__A4 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__B1 (.I(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__A3 (.I(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A2 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__A2 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__A3 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__A4 (.I(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__A2 (.I(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A2 (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A1 (.I(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A2 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A3 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A2 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A4 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A1 (.I(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A2 (.I(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A4 (.I(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__B1 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A2 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A2 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A1 (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A2 (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A1 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A1 (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A2 (.I(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A2 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__A2 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A2 (.I(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__A2 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__A2 (.I(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A2 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__A1 (.I(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__A1 (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A2 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A2 (.I(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__A1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__A2 (.I(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__C (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A2 (.I(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A2 (.I(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A2 (.I(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__A2 (.I(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__A2 (.I(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A2 (.I(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A2 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__A2 (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A1 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A2 (.I(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A2 (.I(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__B1 (.I(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__B2 (.I(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A3 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A2 (.I(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__A1 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__A2 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A3 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A1 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__A2 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__B1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__C1 (.I(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__C2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__A2 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__B1 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__B2 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__B1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__B2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A2 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A1 (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__A2 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A2 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A1 (.I(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A2 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__B1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__B2 (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A1 (.I(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__B1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A1 (.I(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__I (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__A1 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__A2 (.I(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__B2 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A2 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__B1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__B2 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__A1 (.I(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__A1 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__A2 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__B1 (.I(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__B2 (.I(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A2 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A1 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A2 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__B1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A2 (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A1 (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__A3 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A3 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__B (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A2 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A1 (.I(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__B2 (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A2 (.I(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A1 (.I(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A1 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A1 (.I(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A2 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__B1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__B2 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__A1 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__C (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__B1 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__B2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A1 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__A2 (.I(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A1 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__C (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A2 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__B (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A1 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__B (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__I (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A2 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A1 (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__I (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__I (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__I (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A1 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A2 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A1 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A2 (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__I (.I(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A2 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A3 (.I(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A1 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__A3 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__B1 (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__B (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A1 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A2 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__I (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__I (.I(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__I (.I(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A1 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A1 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A1 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__B2 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A1 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__C (.I(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__I (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A1 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__B (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A2 (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A1 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__B (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A2 (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A1 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A2 (.I(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A1 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A1 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A2 (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__C (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A1 (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__B (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A1 (.I(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A1 (.I(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__C (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A1 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__B2 (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__B (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__I (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__B2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__B (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__B2 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__C (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__C (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__I (.I(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A1 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__A2 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__B2 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A1 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A3 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A1 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A1 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A2 (.I(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A1 (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A1 (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__C (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__B2 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__B2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__C (.I(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__B2 (.I(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__B2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A1 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__I (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__C (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__I (.I(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__I0 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__I0 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__I (.I(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__I0 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__I0 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A1 (.I(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A3 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A1 (.I(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A1 (.I(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A2 (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__B (.I(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__I (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A1 (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__B (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__B (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A1 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__I (.I(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A1 (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__A1 (.I(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__B (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__B (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A1 (.I(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__B (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__I (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A1 (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__C (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A1 (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__C (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A1 (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__C (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A1 (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__I (.I(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__A1 (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A1 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__C (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A2 (.I(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A2 (.I(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A3 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A4 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A1 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A3 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__I (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A2 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__I (.I(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__I (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A3 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__I (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__B (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__C (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__I (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__A1 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__B2 (.I(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__I (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__B2 (.I(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__I (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A1 (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__I (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__I (.I(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__I (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__I (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__I (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__I (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__I (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__B2 (.I(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__I (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__B2 (.I(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__A2 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A1 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__I (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A2 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A1 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__A2 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A2 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A2 (.I(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__I (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__I0 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__A1 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A1 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A2 (.I(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A2 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A4 (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A3 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__A1 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__A3 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__B (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__A2 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A2 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A2 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__A2 (.I(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__I (.I(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A2 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A1 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__B2 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A1 (.I(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A3 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A1 (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A2 (.I(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A1 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A1 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__A1 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__A2 (.I(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__B2 (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A1 (.I(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A1 (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A1 (.I(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A1 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A2 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A1 (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__B2 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A1 (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A1 (.I(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A1 (.I(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__A1 (.I(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__B2 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A1 (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A1 (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A2 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__B2 (.I(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__A1 (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A1 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__A1 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__A1 (.I(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__A2 (.I(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__A1 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__B2 (.I(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A2 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__A1 (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__A1 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__A1 (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A1 (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__B1 (.I(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A1 (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A1 (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__A1 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A2 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__B2 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A2 (.I(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A1 (.I(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__I (.I(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A1 (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A3 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__I (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A2 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__B (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__I (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A1 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A2 (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A3 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A2 (.I(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__B1 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__C2 (.I(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__B1 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__C2 (.I(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A2 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__A1 (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A1 (.I(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__B1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__C2 (.I(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__A1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__B1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__I (.I(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A1 (.I(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A1 (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__I (.I(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__B1 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A1 (.I(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11306__B1 (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__B1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__C2 (.I(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A1 (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A1 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__B1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__C2 (.I(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__I (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A2 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A3 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__I (.I(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A2 (.I(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A2 (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__I (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A1 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A1 (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A1 (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__I (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I (.I(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__I (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__A1 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__A1 (.I(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__I (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A2 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__B (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__I (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__I (.I(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__I (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A2 (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A3 (.I(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__A1 (.I(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__B2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__C1 (.I(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__A1 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__B2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__C1 (.I(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A1 (.I(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__B2 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__C1 (.I(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__B2 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__I (.I(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__I (.I(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__I (.I(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__A1 (.I(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__B2 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__A1 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A1 (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__B2 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__A1 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__B2 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__A1 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__B2 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A1 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A1 (.I(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__I (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__A2 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__I (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__I (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A1 (.I(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A2 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__B2 (.I(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A1 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__B2 (.I(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A1 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__B2 (.I(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__A1 (.I(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11390__I (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__I (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__A1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A1 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A1 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__A1 (.I(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A1 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A2 (.I(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__A1 (.I(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__B1 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A2 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__I (.I(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__A1 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A3 (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__A2 (.I(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A1 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A1 (.I(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__B1 (.I(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A1 (.I(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11424__B2 (.I(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A1 (.I(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__B1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__A1 (.I(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__B2 (.I(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A1 (.I(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__B1 (.I(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A1 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__A1 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__B2 (.I(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__I (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11439__A1 (.I(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__A1 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A1 (.I(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__I (.I(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__A1 (.I(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__B2 (.I(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__A1 (.I(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A1 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__C (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__A1 (.I(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__A1 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__B2 (.I(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__C (.I(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__A1 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__A1 (.I(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__B2 (.I(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A1 (.I(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__B1 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__A1 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__A1 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__A4 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__S (.I(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__I0 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__S (.I(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__S (.I(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__I0 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__S (.I(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__S (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__S (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__S (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__I1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__S (.I(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__S (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__S (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__S (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__S (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__I (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11491__S (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__S (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__S (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__S (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__CLK (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__CLK (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__CLK (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11723__CLK (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11886__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11895__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11951__CLK (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__D (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11954__D (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__D (.I(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11956__D (.I(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__D (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11958__D (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11965__D (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__D (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__D (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__D (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__CLK (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__CLK (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12124__I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12125__I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12126__I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12127__I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12131__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_122_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_124_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_128_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_129_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_130_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_131_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_132_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_134_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_135_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_136_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_137_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_138_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_139_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_140_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_141_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_142_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_143_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_144_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_145_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_146_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_147_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_148_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_150_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_151_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_152_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_153_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_154_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_155_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_156_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_157_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_158_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_159_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_160_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_161_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_162_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_163_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_164_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_165_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout258_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout259_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold107_I (.I(wbs_cyc_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold108_I (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold109_I (.I(wbs_dat_i[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold10_I (.I(wbs_dat_i[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold110_I (.I(wbs_dat_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold111_I (.I(wbs_dat_i[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold112_I (.I(wbs_dat_i[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold113_I (.I(wbs_adr_i[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold114_I (.I(wbs_dat_i[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold115_I (.I(wbs_dat_i[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold116_I (.I(wbs_dat_i[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold117_I (.I(wbs_dat_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold118_I (.I(wbs_dat_i[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold119_I (.I(wbs_dat_i[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold11_I (.I(wbs_dat_i[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold120_I (.I(wbs_dat_i[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold121_I (.I(wbs_dat_i[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold122_I (.I(wbs_dat_i[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold123_I (.I(wbs_adr_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold124_I (.I(wbs_dat_i[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold12_I (.I(wbs_dat_i[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold13_I (.I(wbs_dat_i[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold14_I (.I(wbs_dat_i[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold15_I (.I(wbs_dat_i[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold16_I (.I(wbs_dat_i[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold18_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold1_I (.I(wbs_dat_i[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold22_I (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold26_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold2_I (.I(wbs_dat_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold30_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold34_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold3_I (.I(wbs_dat_i[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold48_I (.I(wbs_dat_i[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold4_I (.I(wbs_dat_i[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold5_I (.I(wbs_adr_i[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold65_I (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold67_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold73_I (.I(wbs_dat_i[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold75_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold78_I (.I(wbs_adr_i[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold7_I (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold86_I (.I(wbs_dat_i[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold87_I (.I(wbs_dat_i[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold89_I (.I(wbs_dat_i[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold8_I (.I(wbs_dat_i[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_hold9_I (.I(wbs_dat_i[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(bus_in_serial_ports[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(bus_in_serial_ports[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(bus_in_serial_ports[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(bus_in_serial_ports[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(bus_in_serial_ports[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(bus_in_serial_ports[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(bus_in_serial_ports[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(bus_in_sid[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(bus_in_sid[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(bus_in_sid[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(bus_in_gpios[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(bus_in_sid[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(bus_in_sid[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(bus_in_sid[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(bus_in_sid[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(bus_in_sid[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(bus_in_timers[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(bus_in_timers[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(bus_in_timers[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(bus_in_timers[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(bus_in_timers[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(bus_in_gpios[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(bus_in_timers[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(bus_in_timers[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(bus_in_timers[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(bus_in_gpios[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(irqs[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(irqs[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(irqs[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(irqs[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(irqs[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(irqs[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(irqs[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(bus_in_gpios[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(rom_bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(rom_bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(rom_bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(rom_bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(rom_bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(rom_bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(rom_bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(rom_bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(bus_in_gpios[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_in_gpios[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_in_gpios[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_in_gpios[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input96_I (.I(wbs_stb_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input97_I (.I(wbs_we_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(bus_in_serial_ports[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_max_cap260_I (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output133_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output134_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output147_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output172_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output173_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output177_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output178_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output188_I (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output192_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output198_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output200_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output211_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output213_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output214_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output225_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output245_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output246_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output248_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output249_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer10_I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer12_I (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer13_I (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer1_I (.I(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer2_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer3_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer6_I (.I(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer7_I (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_128_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_168_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_169_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_991 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_615 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05721_ (.I(\as2650.debug_psl[4] ),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05722_ (.I(_00579_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05723_ (.I(_00580_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05724_ (.I(_00581_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05725_ (.I0(\as2650.regs[1][7] ),
    .I1(\as2650.regs[5][7] ),
    .S(_00582_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05726_ (.I(_00583_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05727_ (.I(_00584_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05728_ (.I(_00585_),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05729_ (.I(_00579_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05730_ (.I(_00586_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05731_ (.I0(\as2650.regs[1][6] ),
    .I1(\as2650.regs[5][6] ),
    .S(_00587_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05732_ (.I(_00588_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05733_ (.I(_00589_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05734_ (.I(_00590_),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05735_ (.I(_00587_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05736_ (.I(\as2650.regs[1][5] ),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05737_ (.A1(_00582_),
    .A2(\as2650.regs[5][5] ),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05738_ (.A1(_00591_),
    .A2(_00592_),
    .B(_00593_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05739_ (.I(_00594_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05740_ (.I(_00595_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05741_ (.I(_00596_),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05742_ (.I(_00591_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05743_ (.I(\as2650.regs[1][4] ),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05744_ (.A1(_00591_),
    .A2(\as2650.regs[5][4] ),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05745_ (.A1(_00597_),
    .A2(_00598_),
    .B(_00599_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05746_ (.I(_00600_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05747_ (.I(_00601_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05748_ (.I(_00602_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05749_ (.I(_00603_),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05750_ (.I(\as2650.regs[1][3] ),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05751_ (.A1(_00591_),
    .A2(\as2650.regs[5][3] ),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05752_ (.A1(_00597_),
    .A2(_00604_),
    .B(_00605_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05753_ (.I(_00606_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05754_ (.I(_00607_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05755_ (.I(_00608_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05756_ (.I(_00609_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05757_ (.I(_00610_),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05758_ (.I0(\as2650.regs[1][2] ),
    .I1(\as2650.regs[5][2] ),
    .S(_00580_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05759_ (.I(_00611_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05760_ (.I(_00612_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05761_ (.I(_00613_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05762_ (.I(_00614_),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05763_ (.I0(\as2650.regs[1][1] ),
    .I1(\as2650.regs[5][1] ),
    .S(_00580_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05764_ (.I(_00615_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05765_ (.I(_00616_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05766_ (.I(_00617_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05767_ (.I(_00618_),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05768_ (.I(\as2650.debug_psl[4] ),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05769_ (.I(_00619_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05770_ (.I0(\as2650.regs[1][0] ),
    .I1(\as2650.regs[5][0] ),
    .S(_00620_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05771_ (.I(_00621_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05772_ (.I(_00622_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05773_ (.I(_00623_),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05774_ (.I(\as2650.debug_psl[4] ),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05775_ (.I(_00624_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05776_ (.I(_00625_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05777_ (.A1(_00582_),
    .A2(\as2650.regs[0][7] ),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05778_ (.A1(_00626_),
    .A2(\as2650.regs[4][7] ),
    .B(_00627_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05779_ (.I(_00628_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05780_ (.I(_00629_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05781_ (.I(_00630_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05782_ (.I(_00631_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05783_ (.I(_00632_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05784_ (.I(_00633_),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05785_ (.I(_00579_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05786_ (.I(\as2650.regs[4][6] ),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05787_ (.A1(_00634_),
    .A2(_00635_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05788_ (.A1(_00586_),
    .A2(\as2650.regs[0][6] ),
    .B(_00636_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05789_ (.I(_00637_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05790_ (.I(_00638_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05791_ (.I(_00639_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05792_ (.I(_00640_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05793_ (.I(_00641_),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05794_ (.I(_00642_),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05795_ (.I(\as2650.regs[4][5] ),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05796_ (.A1(_00619_),
    .A2(_00643_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05797_ (.A1(_00580_),
    .A2(\as2650.regs[0][5] ),
    .B(_00644_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05798_ (.I(_00645_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05799_ (.I(_00646_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05800_ (.I(_00647_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05801_ (.I(_00648_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05802_ (.I(_00649_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05803_ (.I(_00650_),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05804_ (.I(\as2650.regs[4][4] ),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05805_ (.A1(_00579_),
    .A2(_00651_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05806_ (.A1(_00619_),
    .A2(\as2650.regs[0][4] ),
    .B(_00652_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05807_ (.I(_00653_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05808_ (.I(_00654_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05809_ (.I(_00655_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05810_ (.I(_00656_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05811_ (.I(_00657_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05812_ (.I(_00658_),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05813_ (.I(\as2650.cycle[3] ),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05814_ (.I(_00659_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05815_ (.I(\as2650.cycle[1] ),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05816_ (.I(_00661_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05817_ (.I(_00662_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05818_ (.I(_00663_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05819_ (.I(\as2650.cycle[2] ),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05820_ (.A1(_00664_),
    .A2(_00665_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05821_ (.A1(_00660_),
    .A2(_00666_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05822_ (.I(_00667_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05823_ (.I(_00668_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05824_ (.A1(\as2650.cycle[2] ),
    .A2(\as2650.cycle[3] ),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05825_ (.I(\as2650.cycle[0] ),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05826_ (.A1(_00671_),
    .A2(_00661_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05827_ (.A1(_00670_),
    .A2(_00672_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05828_ (.I(_00673_),
    .Z(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05829_ (.I(\as2650.relative_cyc ),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05830_ (.I(_00665_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05831_ (.I(\as2650.indirect_cyc ),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05832_ (.A1(_00661_),
    .A2(_00676_),
    .A3(_00660_),
    .B(_00677_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05833_ (.I(_00678_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05834_ (.A1(_00675_),
    .A2(_00679_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _05835_ (.A1(_00674_),
    .A2(_00680_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05836_ (.I(_00671_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05837_ (.A1(_00665_),
    .A2(_00659_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05838_ (.A1(_00682_),
    .A2(_00662_),
    .A3(_00683_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05839_ (.A1(\as2650.indexed_cyc[1] ),
    .A2(\as2650.indexed_cyc[0] ),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05840_ (.A1(\as2650.wb_hidden_rom_enable ),
    .A2(\as2650.cpu_hidden_rom_enable ),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05841_ (.I(_00686_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05842_ (.I(\as2650.wb_hidden_rom_enable ),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05843_ (.I(_00688_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05844_ (.I(\as2650.cpu_hidden_rom_enable ),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05845_ (.A1(_00689_),
    .A2(_00690_),
    .A3(net57),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__or4_4 _05846_ (.A1(\as2650.cycle[0] ),
    .A2(\as2650.cycle[1] ),
    .A3(\as2650.cycle[2] ),
    .A4(\as2650.cycle[3] ),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05847_ (.I(_00692_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05848_ (.I(_00693_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05849_ (.A1(net36),
    .A2(_00687_),
    .B(_00691_),
    .C(_00694_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05850_ (.A1(_00671_),
    .A2(_00661_),
    .A3(net319),
    .A4(net318),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05851_ (.I(_00696_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05852_ (.A1(\as2650.insin[7] ),
    .A2(_00697_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05853_ (.I(_00693_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05854_ (.A1(\as2650.insin[6] ),
    .A2(_00699_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05855_ (.I(net56),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05856_ (.I(_00686_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05857_ (.I(_00702_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05858_ (.I(_00689_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05859_ (.I(_00690_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05860_ (.A1(_00704_),
    .A2(_00705_),
    .B(net35),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05861_ (.A1(_00701_),
    .A2(_00703_),
    .B(_00706_),
    .C(_00694_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05862_ (.A1(_00695_),
    .A2(_00698_),
    .A3(_00700_),
    .A4(_00707_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05863_ (.A1(\as2650.insin[4] ),
    .A2(_00699_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05864_ (.I(net54),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05865_ (.I(_00703_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05866_ (.I(_00689_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05867_ (.I(_00690_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05868_ (.A1(_00712_),
    .A2(_00713_),
    .B(net42),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05869_ (.A1(_00710_),
    .A2(_00711_),
    .B(_00714_),
    .C(_00699_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05870_ (.A1(\as2650.insin[5] ),
    .A2(_00699_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _05871_ (.I(net55),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05872_ (.A1(_00704_),
    .A2(_00713_),
    .B(net34),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05873_ (.A1(_00717_),
    .A2(_00703_),
    .B(_00718_),
    .C(_00694_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05874_ (.A1(_00709_),
    .A2(_00715_),
    .A3(_00716_),
    .A4(_00719_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05875_ (.I(_00694_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05876_ (.A1(\as2650.insin[7] ),
    .A2(_00721_),
    .Z(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05877_ (.I(net57),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05878_ (.A1(_00712_),
    .A2(_00713_),
    .B(net36),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05879_ (.I(_00693_),
    .Z(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05880_ (.A1(_00723_),
    .A2(_00711_),
    .B(_00724_),
    .C(_00725_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _05881_ (.A1(_00704_),
    .A2(_00705_),
    .A3(net56),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05882_ (.A1(net35),
    .A2(_00687_),
    .B(_00727_),
    .C(_00725_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05883_ (.A1(\as2650.insin[6] ),
    .A2(_00697_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05884_ (.A1(_00722_),
    .A2(_00726_),
    .A3(_00728_),
    .A4(_00729_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05885_ (.I(\as2650.extend ),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05886_ (.A1(_00708_),
    .A2(_00720_),
    .A3(_00730_),
    .B(_00731_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05887_ (.I(\as2650.indirect_cyc ),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _05888_ (.A1(_00689_),
    .A2(_00705_),
    .A3(net53),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05889_ (.A1(net41),
    .A2(_00687_),
    .B(_00734_),
    .C(_00725_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05890_ (.A1(\as2650.insin[3] ),
    .A2(_00697_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05891_ (.A1(_00735_),
    .A2(_00736_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05892_ (.I0(net40),
    .I1(net52),
    .S(_00711_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05893_ (.I(_00696_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05894_ (.A1(\as2650.insin[2] ),
    .A2(_00739_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05895_ (.A1(_00721_),
    .A2(_00738_),
    .B(_00740_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05896_ (.A1(_00733_),
    .A2(_00737_),
    .A3(_00741_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05897_ (.I(_00687_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _05898_ (.A1(_00704_),
    .A2(_00705_),
    .A3(net54),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05899_ (.A1(net42),
    .A2(_00743_),
    .B(_00744_),
    .C(_00725_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05900_ (.A1(\as2650.insin[4] ),
    .A2(_00697_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05901_ (.A1(_00745_),
    .A2(_00746_),
    .A3(_00735_),
    .A4(_00736_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05902_ (.I(\as2650.instruction_args_latch[13] ),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05903_ (.A1(_00748_),
    .A2(\as2650.instruction_args_latch[14] ),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05904_ (.I(\as2650.extend ),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05905_ (.A1(_00747_),
    .A2(_00749_),
    .B(_00750_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05906_ (.A1(_00732_),
    .A2(_00742_),
    .A3(_00751_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05907_ (.A1(_00684_),
    .A2(_00685_),
    .B(_00752_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05908_ (.A1(_00681_),
    .A2(_00753_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05909_ (.I(_00754_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05910_ (.I(\as2650.instruction_args_latch[14] ),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05911_ (.I(\as2650.indexed_cyc[1] ),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05912_ (.A1(\as2650.indexed_cyc[0] ),
    .A2(_00756_),
    .B(_00757_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05913_ (.A1(\as2650.extend ),
    .A2(_00758_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05914_ (.I(\as2650.instruction_args_latch[13] ),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05915_ (.I(\as2650.indexed_cyc[0] ),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _05916_ (.A1(\as2650.indexed_cyc[1] ),
    .A2(_00760_),
    .B(_00761_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05917_ (.A1(_00759_),
    .A2(_00762_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05918_ (.I(_00763_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05919_ (.A1(_00688_),
    .A2(net50),
    .A3(\as2650.cpu_hidden_rom_enable ),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _05920_ (.I(_00692_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05921_ (.A1(net38),
    .A2(_00686_),
    .B(_00765_),
    .C(_00766_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05922_ (.A1(\as2650.insin[0] ),
    .A2(_00696_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05923_ (.A1(net310),
    .A2(_00768_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05924_ (.I(_00769_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05925_ (.I(_00770_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05926_ (.A1(\as2650.insin[0] ),
    .A2(_00693_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05927_ (.I(_00772_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05928_ (.I(net50),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05929_ (.A1(_00688_),
    .A2(_00690_),
    .B(net38),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05930_ (.A1(_00774_),
    .A2(_00703_),
    .B(_00775_),
    .C(_00766_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05931_ (.I(net304),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05932_ (.A1(_00773_),
    .A2(_00777_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05933_ (.I(_00778_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05934_ (.A1(\as2650.regs[6][7] ),
    .A2(_00779_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05935_ (.A1(\as2650.insin[1] ),
    .A2(_00766_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05936_ (.I(_00781_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05937_ (.I(net51),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05938_ (.A1(_00688_),
    .A2(\as2650.cpu_hidden_rom_enable ),
    .B(net39),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05939_ (.A1(_00783_),
    .A2(_00702_),
    .B(_00784_),
    .C(_00766_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05940_ (.I(net307),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05941_ (.A1(_00782_),
    .A2(_00786_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05942_ (.I(_00787_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05943_ (.I(_00788_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05944_ (.A1(\as2650.regs[7][7] ),
    .A2(_00771_),
    .B(_00780_),
    .C(_00789_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05945_ (.I(_00767_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05946_ (.A1(_00782_),
    .A2(_00786_),
    .A3(_00791_),
    .A4(_00768_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05947_ (.I(_00792_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05948_ (.I(_00793_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05949_ (.A1(_00782_),
    .A2(_00786_),
    .A3(_00772_),
    .A4(net305),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05950_ (.I(_00795_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05951_ (.I(_00796_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05952_ (.I(_00586_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05953_ (.A1(\as2650.regs[5][7] ),
    .A2(_00794_),
    .B1(_00797_),
    .B2(\as2650.regs[4][7] ),
    .C(_00798_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05954_ (.I(_00778_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05955_ (.A1(\as2650.regs[2][7] ),
    .A2(_00800_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05956_ (.I(_00788_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05957_ (.A1(\as2650.regs[3][7] ),
    .A2(_00771_),
    .B(_00801_),
    .C(_00802_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05958_ (.I(_00793_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05959_ (.I(_00796_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _05960_ (.A1(\as2650.regs[1][7] ),
    .A2(_00804_),
    .B1(_00805_),
    .B2(\as2650.regs[0][7] ),
    .C(_00626_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05961_ (.A1(_00790_),
    .A2(_00799_),
    .B1(_00803_),
    .B2(_00806_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05962_ (.I(_00807_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _05963_ (.A1(_00782_),
    .A2(_00786_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05964_ (.I(_00809_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05965_ (.I(_00810_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05966_ (.I0(\as2650.regs[7][6] ),
    .I1(\as2650.regs[6][6] ),
    .S(_00800_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _05967_ (.I(_00795_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05968_ (.A1(_00635_),
    .A2(_00813_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05969_ (.I(\as2650.regs[5][6] ),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05970_ (.I(_00792_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05971_ (.A1(_00815_),
    .A2(_00816_),
    .B(_00620_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05972_ (.A1(_00811_),
    .A2(_00812_),
    .B(_00814_),
    .C(_00817_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05973_ (.I0(\as2650.regs[3][6] ),
    .I1(\as2650.regs[2][6] ),
    .S(_00800_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05974_ (.I(\as2650.regs[0][6] ),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05975_ (.I(_00791_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05976_ (.I(_00768_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05977_ (.A1(\as2650.regs[1][6] ),
    .A2(_00821_),
    .A3(_00822_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05978_ (.A1(_00820_),
    .A2(_00779_),
    .B(_00823_),
    .C(_00810_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05979_ (.A1(_00811_),
    .A2(_00819_),
    .B(_00824_),
    .C(_00587_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05980_ (.A1(_00818_),
    .A2(_00825_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05981_ (.I(\as2650.regs[7][5] ),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05982_ (.I(_00769_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05983_ (.I(_00773_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05984_ (.I(_00777_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05985_ (.A1(\as2650.regs[6][5] ),
    .A2(_00829_),
    .A3(_00830_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05986_ (.I(_00787_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05987_ (.A1(_00827_),
    .A2(_00828_),
    .B(_00831_),
    .C(_00832_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05988_ (.I(\as2650.regs[5][5] ),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05989_ (.A1(_00834_),
    .A2(_00816_),
    .B1(_00813_),
    .B2(_00643_),
    .C(_00620_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05990_ (.I(\as2650.regs[2][5] ),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05991_ (.A1(\as2650.regs[3][5] ),
    .A2(_00791_),
    .A3(_00822_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05992_ (.A1(_00836_),
    .A2(_00800_),
    .B(_00837_),
    .C(_00788_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05993_ (.I(\as2650.regs[0][5] ),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05994_ (.I(_00624_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _05995_ (.A1(_00592_),
    .A2(_00816_),
    .B1(_00813_),
    .B2(_00839_),
    .C(_00840_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05996_ (.A1(_00833_),
    .A2(_00835_),
    .B1(_00838_),
    .B2(_00841_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05997_ (.I(_00842_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05998_ (.I(\as2650.regs[7][4] ),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05999_ (.I(_00769_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06000_ (.I(_00773_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06001_ (.I(_00777_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06002_ (.A1(\as2650.regs[6][4] ),
    .A2(_00846_),
    .A3(_00847_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06003_ (.A1(_00844_),
    .A2(_00845_),
    .B(_00848_),
    .C(_00832_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06004_ (.I(\as2650.regs[5][4] ),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06005_ (.A1(_00850_),
    .A2(_00793_),
    .B1(_00796_),
    .B2(_00651_),
    .C(_00586_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06006_ (.I(\as2650.regs[2][4] ),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06007_ (.A1(\as2650.regs[3][4] ),
    .A2(_00791_),
    .A3(_00822_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06008_ (.A1(_00852_),
    .A2(_00778_),
    .B(_00853_),
    .C(_00788_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06009_ (.I(\as2650.regs[0][4] ),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06010_ (.A1(_00598_),
    .A2(_00793_),
    .B1(_00796_),
    .B2(_00855_),
    .C(_00840_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06011_ (.A1(_00849_),
    .A2(_00851_),
    .B1(_00854_),
    .B2(_00856_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06012_ (.I(_00857_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06013_ (.I(\as2650.regs[6][1] ),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06014_ (.I(_00772_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06015_ (.I(net306),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06016_ (.A1(_00860_),
    .A2(_00861_),
    .B(\as2650.regs[7][1] ),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06017_ (.I(_00809_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06018_ (.A1(_00859_),
    .A2(_00845_),
    .B(_00862_),
    .C(_00863_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06019_ (.I(\as2650.regs[5][1] ),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06020_ (.A1(_00781_),
    .A2(net307),
    .A3(net313),
    .A4(_00768_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06021_ (.I(_00866_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06022_ (.A1(_00781_),
    .A2(net307),
    .A3(_00772_),
    .A4(net316),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06023_ (.I(_00868_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06024_ (.I(\as2650.regs[4][1] ),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06025_ (.A1(_00865_),
    .A2(_00867_),
    .B1(_00869_),
    .B2(_00870_),
    .C(_00625_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06026_ (.I(\as2650.regs[2][1] ),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06027_ (.A1(_00846_),
    .A2(_00847_),
    .B(\as2650.regs[3][1] ),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06028_ (.A1(_00872_),
    .A2(_00845_),
    .B(_00873_),
    .C(_00863_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06029_ (.I(\as2650.regs[1][1] ),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06030_ (.I(\as2650.regs[0][1] ),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06031_ (.A1(_00875_),
    .A2(_00867_),
    .B1(_00869_),
    .B2(_00876_),
    .C(_00634_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06032_ (.A1(_00864_),
    .A2(_00871_),
    .B1(_00874_),
    .B2(_00877_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06033_ (.I(\as2650.regs[6][0] ),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06034_ (.A1(_00846_),
    .A2(_00847_),
    .B(\as2650.regs[7][0] ),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06035_ (.A1(_00879_),
    .A2(_00845_),
    .B(_00880_),
    .C(_00810_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06036_ (.I(\as2650.regs[5][0] ),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06037_ (.I(\as2650.regs[4][0] ),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06038_ (.A1(_00882_),
    .A2(_00867_),
    .B1(_00869_),
    .B2(_00883_),
    .C(_00625_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06039_ (.I(\as2650.regs[2][0] ),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06040_ (.A1(_00846_),
    .A2(_00847_),
    .B(\as2650.regs[3][0] ),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06041_ (.A1(_00885_),
    .A2(_00828_),
    .B(_00886_),
    .C(_00810_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06042_ (.I(\as2650.regs[1][0] ),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06043_ (.I(_00866_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06044_ (.I(_00889_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06045_ (.I(_00868_),
    .Z(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06046_ (.I(_00891_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06047_ (.I(\as2650.regs[0][0] ),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06048_ (.A1(_00888_),
    .A2(_00890_),
    .B1(_00892_),
    .B2(_00893_),
    .C(_00634_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06049_ (.A1(_00881_),
    .A2(_00884_),
    .B1(_00887_),
    .B2(_00894_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06050_ (.I(\as2650.regs[6][3] ),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06051_ (.A1(_00860_),
    .A2(_00861_),
    .B(\as2650.regs[7][3] ),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06052_ (.A1(_00896_),
    .A2(_00770_),
    .B(_00897_),
    .C(_00863_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06053_ (.I(\as2650.regs[5][3] ),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06054_ (.I(\as2650.regs[4][3] ),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06055_ (.A1(_00899_),
    .A2(net317),
    .B1(net311),
    .B2(_00900_),
    .C(_00625_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06056_ (.I(\as2650.regs[2][3] ),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06057_ (.A1(_00860_),
    .A2(_00861_),
    .B(\as2650.regs[3][3] ),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06058_ (.A1(_00902_),
    .A2(_00770_),
    .B(_00903_),
    .C(_00863_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06059_ (.I(\as2650.regs[0][3] ),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06060_ (.A1(_00604_),
    .A2(_00867_),
    .B1(_00869_),
    .B2(_00905_),
    .C(_00634_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06061_ (.A1(_00898_),
    .A2(_00901_),
    .B1(_00904_),
    .B2(_00906_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06062_ (.I(\as2650.regs[6][2] ),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06063_ (.A1(_00860_),
    .A2(_00861_),
    .B(\as2650.regs[7][2] ),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06064_ (.A1(_00908_),
    .A2(_00770_),
    .B(_00909_),
    .C(_00809_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06065_ (.I(\as2650.regs[5][2] ),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06066_ (.I(\as2650.regs[4][2] ),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06067_ (.A1(_00911_),
    .A2(net317),
    .B1(net312),
    .B2(_00912_),
    .C(_00624_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06068_ (.I(\as2650.regs[2][2] ),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06069_ (.A1(_00773_),
    .A2(_00777_),
    .B(\as2650.regs[3][2] ),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06070_ (.A1(_00914_),
    .A2(_00769_),
    .B(_00915_),
    .C(_00809_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06071_ (.I(\as2650.regs[1][2] ),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06072_ (.I(\as2650.regs[0][2] ),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06073_ (.A1(_00917_),
    .A2(net317),
    .B1(net311),
    .B2(_00918_),
    .C(_00619_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06074_ (.A1(_00910_),
    .A2(_00913_),
    .B1(_00916_),
    .B2(_00919_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06075_ (.A1(_00878_),
    .A2(_00895_),
    .A3(_00907_),
    .A4(_00920_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06076_ (.A1(_00826_),
    .A2(_00843_),
    .A3(_00858_),
    .A4(_00921_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06077_ (.A1(_00808_),
    .A2(_00922_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06078_ (.A1(_00764_),
    .A2(_00923_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06079_ (.A1(\as2650.extend ),
    .A2(_00762_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06080_ (.A1(_00758_),
    .A2(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06081_ (.I(_00926_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06082_ (.I(_00807_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06083_ (.A1(_00818_),
    .A2(_00825_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06084_ (.I(_00920_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06085_ (.A1(_00878_),
    .A2(_00895_),
    .A3(_00907_),
    .A4(_00930_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06086_ (.A1(_00842_),
    .A2(_00858_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06087_ (.A1(_00929_),
    .A2(_00931_),
    .A3(_00932_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06088_ (.A1(_00928_),
    .A2(_00933_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06089_ (.A1(_00808_),
    .A2(_00927_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06090_ (.A1(_00927_),
    .A2(_00934_),
    .B(_00935_),
    .C(_00764_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__and3_4 _06091_ (.A1(_00755_),
    .A2(_00924_),
    .A3(_00936_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _06092_ (.A1(_00675_),
    .A2(_00733_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06093_ (.I(_00938_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06094_ (.I(_00939_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06095_ (.I(_00670_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06096_ (.A1(_00675_),
    .A2(_00941_),
    .A3(_00674_),
    .A4(_00679_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06097_ (.I(net264),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06098_ (.A1(\as2650.indirect_target[7] ),
    .A2(_00940_),
    .B1(_00943_),
    .B2(\as2650.PC[7] ),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06099_ (.A1(\as2650.indirect_target[6] ),
    .A2(_00940_),
    .B1(_00943_),
    .B2(\as2650.PC[6] ),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06100_ (.A1(\as2650.indirect_target[5] ),
    .A2(_00939_),
    .B1(_00943_),
    .B2(\as2650.PC[5] ),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06101_ (.I(_00946_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06102_ (.A1(\as2650.indirect_target[4] ),
    .A2(_00939_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06103_ (.A1(\as2650.PC[4] ),
    .A2(net264),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06104_ (.A1(_00948_),
    .A2(_00949_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06105_ (.I(\as2650.PC[3] ),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06106_ (.A1(\as2650.relative_cyc ),
    .A2(_00941_),
    .A3(_00673_),
    .A4(_00678_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06107_ (.I(_00952_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06108_ (.A1(\as2650.indirect_target[3] ),
    .A2(_00939_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06109_ (.A1(_00951_),
    .A2(_00953_),
    .B(_00954_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06110_ (.A1(\as2650.indirect_target[1] ),
    .A2(_00938_),
    .B1(_00942_),
    .B2(\as2650.PC[1] ),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06111_ (.I(\as2650.PC[0] ),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06112_ (.A1(\as2650.indirect_target[0] ),
    .A2(_00938_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06113_ (.I0(_00957_),
    .I1(_00958_),
    .S(_00952_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06114_ (.A1(_00671_),
    .A2(_00663_),
    .A3(_00941_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06115_ (.A1(_00680_),
    .A2(_00960_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06116_ (.A1(\as2650.indirect_target[2] ),
    .A2(_00938_),
    .B1(net264),
    .B2(\as2650.PC[2] ),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06117_ (.A1(_00956_),
    .A2(_00959_),
    .A3(_00961_),
    .A4(_00962_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06118_ (.A1(_00947_),
    .A2(_00950_),
    .A3(_00955_),
    .A4(_00963_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06119_ (.A1(_00945_),
    .A2(_00964_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06120_ (.A1(_00944_),
    .A2(_00965_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06121_ (.I(_00684_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06122_ (.A1(_00944_),
    .A2(_00965_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06123_ (.A1(_00967_),
    .A2(_00968_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06124_ (.I(_00674_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06125_ (.I(_00970_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06126_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_00971_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06127_ (.A1(_00966_),
    .A2(_00969_),
    .B(_00972_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06128_ (.A1(_00973_),
    .A2(_00937_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06129_ (.A1(_00681_),
    .A2(_00753_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06130_ (.I(_00975_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06131_ (.I(_00926_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06132_ (.I(_00895_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06133_ (.A1(_00878_),
    .A2(_00978_),
    .A3(_00907_),
    .A4(_00930_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06134_ (.I(_00857_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06135_ (.A1(_00843_),
    .A2(_00980_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06136_ (.A1(_00979_),
    .A2(_00981_),
    .B(_00826_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06137_ (.I(_00926_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06138_ (.I(_00826_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06139_ (.A1(_00983_),
    .A2(_00984_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06140_ (.A1(_00977_),
    .A2(_00933_),
    .A3(_00982_),
    .B(_00985_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__or3_4 _06141_ (.A1(_00843_),
    .A2(_00858_),
    .A3(_00921_),
    .Z(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06142_ (.A1(_00929_),
    .A2(_00987_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06143_ (.A1(_00759_),
    .A2(_00762_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _06144_ (.I0(_00986_),
    .I1(_00988_),
    .S(_00989_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _06145_ (.A1(_00976_),
    .A2(_00990_),
    .Z(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06146_ (.I(_00970_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06147_ (.A1(_00945_),
    .A2(_00964_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06148_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_00992_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06149_ (.A1(_00992_),
    .A2(_00993_),
    .B(_00994_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06150_ (.A1(_00991_),
    .A2(_00995_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06151_ (.A1(_00879_),
    .A2(_00829_),
    .A3(_00830_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06152_ (.A1(\as2650.regs[7][0] ),
    .A2(_00771_),
    .B(_00997_),
    .C(_00789_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06153_ (.I(\as2650.regs[4][0] ),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06154_ (.A1(\as2650.regs[5][0] ),
    .A2(_00794_),
    .B1(_00797_),
    .B2(_00999_),
    .C(_00798_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06155_ (.I(_00778_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06156_ (.I(\as2650.regs[3][0] ),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06157_ (.I(_00822_),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06158_ (.A1(_01002_),
    .A2(_00821_),
    .A3(_01003_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06159_ (.A1(\as2650.regs[2][0] ),
    .A2(_01001_),
    .B(_01004_),
    .C(_00802_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06160_ (.I(\as2650.regs[0][0] ),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06161_ (.A1(\as2650.regs[1][0] ),
    .A2(_00794_),
    .B1(_00797_),
    .B2(_01006_),
    .C(_00626_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06162_ (.A1(_00998_),
    .A2(_01000_),
    .B1(_01005_),
    .B2(_01007_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06163_ (.I(_01008_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06164_ (.I(_00763_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06165_ (.A1(_01010_),
    .A2(_00983_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06166_ (.A1(_01009_),
    .A2(_01011_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06167_ (.I(_00674_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06168_ (.A1(_00959_),
    .A2(_00961_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06169_ (.A1(_00959_),
    .A2(_00961_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06170_ (.A1(\as2650.instruction_args_latch[0] ),
    .A2(_00970_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06171_ (.A1(_01013_),
    .A2(_01014_),
    .A3(_01015_),
    .B(_01016_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06172_ (.A1(_00755_),
    .A2(_01012_),
    .A3(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06173_ (.A1(_00859_),
    .A2(_00829_),
    .A3(_00830_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06174_ (.A1(\as2650.regs[7][1] ),
    .A2(_00828_),
    .B(_01019_),
    .C(_00832_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06175_ (.A1(\as2650.regs[5][1] ),
    .A2(_00804_),
    .B1(_00805_),
    .B2(\as2650.regs[4][1] ),
    .C(_00581_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06176_ (.I(\as2650.regs[3][1] ),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06177_ (.A1(_01022_),
    .A2(_00821_),
    .A3(_01003_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06178_ (.A1(\as2650.regs[2][1] ),
    .A2(_00779_),
    .B(_01023_),
    .C(_00832_),
    .ZN(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06179_ (.I(\as2650.regs[0][1] ),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06180_ (.A1(\as2650.regs[1][1] ),
    .A2(_00816_),
    .B1(_00813_),
    .B2(_01025_),
    .C(_00840_),
    .ZN(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06181_ (.A1(_01020_),
    .A2(_01021_),
    .B1(_01024_),
    .B2(_01026_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06182_ (.A1(_01027_),
    .A2(_00978_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06183_ (.A1(_00758_),
    .A2(_00925_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06184_ (.A1(_01029_),
    .A2(_01009_),
    .B(_00763_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _06185_ (.A1(_01030_),
    .A2(_01028_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06186_ (.A1(_00956_),
    .A2(_01014_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06187_ (.A1(\as2650.instruction_args_latch[1] ),
    .A2(_00970_),
    .ZN(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06188_ (.A1(_00976_),
    .A2(_01031_),
    .B1(_01032_),
    .B2(_00992_),
    .C(_01033_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06189_ (.A1(_01030_),
    .A2(_01028_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06190_ (.A1(_01013_),
    .A2(_01032_),
    .B(_01033_),
    .ZN(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06191_ (.A1(_00755_),
    .A2(_01035_),
    .A3(_01036_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06192_ (.A1(_01018_),
    .A2(_01034_),
    .B(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06193_ (.I(_01010_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06194_ (.A1(_00908_),
    .A2(_00829_),
    .A3(_00830_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06195_ (.A1(\as2650.regs[7][2] ),
    .A2(_00828_),
    .B(_01040_),
    .C(_00802_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06196_ (.A1(\as2650.regs[5][2] ),
    .A2(_00804_),
    .B1(_00805_),
    .B2(\as2650.regs[4][2] ),
    .C(_00798_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06197_ (.I(\as2650.regs[3][2] ),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06198_ (.A1(_01043_),
    .A2(_00821_),
    .A3(_01003_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06199_ (.A1(\as2650.regs[2][2] ),
    .A2(_00779_),
    .B(_01044_),
    .C(_00802_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06200_ (.I(\as2650.regs[0][2] ),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06201_ (.A1(\as2650.regs[1][2] ),
    .A2(_00804_),
    .B1(_00805_),
    .B2(_01046_),
    .C(_00840_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06202_ (.A1(_01041_),
    .A2(_01042_),
    .B1(_01045_),
    .B2(_01047_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06203_ (.A1(_01027_),
    .A2(_01008_),
    .A3(_01048_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06204_ (.I(_01049_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06205_ (.I(_00878_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06206_ (.A1(_01051_),
    .A2(_00978_),
    .B(_00930_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06207_ (.I(_00930_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06208_ (.A1(_00983_),
    .A2(_01053_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06209_ (.A1(_00977_),
    .A2(_01050_),
    .A3(_01052_),
    .B(_01054_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06210_ (.A1(_01027_),
    .A2(_01008_),
    .A3(_01048_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06211_ (.I(_00978_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06212_ (.A1(_01051_),
    .A2(_01057_),
    .B(_01053_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06213_ (.A1(_01056_),
    .A2(_01058_),
    .B(_01010_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06214_ (.A1(_01039_),
    .A2(_01055_),
    .B(_01059_),
    .C(_00975_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06215_ (.A1(_00956_),
    .A2(_00959_),
    .A3(_00961_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06216_ (.A1(_01061_),
    .A2(_00962_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06217_ (.A1(\as2650.instruction_args_latch[2] ),
    .A2(_01013_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06218_ (.A1(_00971_),
    .A2(_01062_),
    .B(_01063_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06219_ (.I(_01064_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06220_ (.A1(_01060_),
    .A2(_01065_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06221_ (.I(_01060_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06222_ (.A1(_01067_),
    .A2(_01064_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06223_ (.A1(_01038_),
    .A2(_01066_),
    .B(_01068_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06224_ (.I(_00907_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06225_ (.I(_00931_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06226_ (.A1(_01070_),
    .A2(_01049_),
    .B(_01071_),
    .C(_01029_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06227_ (.A1(_00983_),
    .A2(_01070_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06228_ (.A1(_01010_),
    .A2(_01072_),
    .A3(_01073_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06229_ (.A1(_00898_),
    .A2(_00901_),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06230_ (.A1(_00904_),
    .A2(_00906_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06231_ (.A1(_01075_),
    .A2(_01076_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06232_ (.A1(_01077_),
    .A2(_01056_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06233_ (.A1(_00764_),
    .A2(_01078_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06234_ (.A1(_01074_),
    .A2(_01079_),
    .B(_00754_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06235_ (.A1(_00955_),
    .A2(_00963_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06236_ (.A1(_00955_),
    .A2(_00963_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06237_ (.A1(_01013_),
    .A2(_01081_),
    .A3(_01082_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06238_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_00971_),
    .B(_01083_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06239_ (.A1(_01080_),
    .A2(_01084_),
    .Z(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06240_ (.A1(_01080_),
    .A2(_01084_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06241_ (.A1(_01069_),
    .A2(_01085_),
    .B(_01086_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06242_ (.A1(_01071_),
    .A2(_00932_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06243_ (.I(_00843_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06244_ (.A1(_00979_),
    .A2(_00980_),
    .B(_01089_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06245_ (.A1(_00977_),
    .A2(_01089_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06246_ (.A1(_00927_),
    .A2(_01088_),
    .A3(_01090_),
    .B(_01091_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06247_ (.I(_00980_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06248_ (.A1(_01093_),
    .A2(_00921_),
    .B(_01089_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06249_ (.A1(_00987_),
    .A2(_01094_),
    .B(_00764_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06250_ (.A1(_01039_),
    .A2(_01092_),
    .B(_01095_),
    .C(_00975_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06251_ (.A1(_00950_),
    .A2(_01081_),
    .B(_00947_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06252_ (.A1(_00967_),
    .A2(_00964_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06253_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_00971_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06254_ (.A1(_01097_),
    .A2(_01098_),
    .B(_01099_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06255_ (.A1(_01096_),
    .A2(_01100_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06256_ (.A1(_01071_),
    .A2(_00980_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06257_ (.A1(_00977_),
    .A2(_01093_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06258_ (.A1(_00927_),
    .A2(_01102_),
    .B(_01103_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06259_ (.A1(_00921_),
    .A2(_00858_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06260_ (.A1(_00989_),
    .A2(_01105_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06261_ (.A1(_01039_),
    .A2(_01104_),
    .B(_01106_),
    .C(_00976_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06262_ (.A1(_00950_),
    .A2(_01081_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06263_ (.I0(\as2650.instruction_args_latch[4] ),
    .I1(_01108_),
    .S(_00967_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06264_ (.A1(_01109_),
    .A2(_01107_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06265_ (.A1(_01110_),
    .A2(_01101_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06266_ (.A1(_00974_),
    .A2(_00996_),
    .A3(_01087_),
    .A4(_01111_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06267_ (.I(_01112_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06268_ (.A1(_01096_),
    .A2(_01100_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06269_ (.A1(_01107_),
    .A2(_01109_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06270_ (.A1(_01096_),
    .A2(_01100_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06271_ (.A1(_01114_),
    .A2(_01115_),
    .B(_01116_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06272_ (.I(_00995_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06273_ (.A1(_00976_),
    .A2(_00990_),
    .A3(_01118_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06274_ (.A1(_00937_),
    .A2(_00973_),
    .B(_01119_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06275_ (.A1(_00937_),
    .A2(_00973_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _06276_ (.A1(_00974_),
    .A2(_00996_),
    .A3(_01117_),
    .B1(_01120_),
    .B2(_01121_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06277_ (.I(_01122_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06278_ (.I(_00992_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06279_ (.I(_01124_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06280_ (.I(_00943_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06281_ (.A1(\as2650.indirect_target[8] ),
    .A2(_00940_),
    .B1(_01126_),
    .B2(\as2650.PC[8] ),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06282_ (.A1(_00944_),
    .A2(_00945_),
    .A3(_00964_),
    .A4(_01127_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06283_ (.I(_00940_),
    .Z(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06284_ (.A1(\as2650.indirect_target[9] ),
    .A2(_01129_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06285_ (.A1(\as2650.PC[9] ),
    .A2(_01126_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06286_ (.A1(_01130_),
    .A2(_01131_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06287_ (.A1(_01128_),
    .A2(_01132_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06288_ (.I(_01133_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06289_ (.A1(\as2650.indirect_target[10] ),
    .A2(_01129_),
    .B1(_01126_),
    .B2(\as2650.PC[10] ),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06290_ (.I(_01135_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06291_ (.I(_01126_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06292_ (.A1(\as2650.indirect_target[11] ),
    .A2(_01129_),
    .B1(_01137_),
    .B2(\as2650.PC[11] ),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06293_ (.A1(_01134_),
    .A2(_01136_),
    .B(_01138_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06294_ (.I(_01124_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06295_ (.A1(_01133_),
    .A2(_01136_),
    .A3(_01138_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06296_ (.A1(_01140_),
    .A2(_01141_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06297_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(_01125_),
    .B1(_01139_),
    .B2(_01142_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06298_ (.A1(_01134_),
    .A2(_01136_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06299_ (.A1(_01134_),
    .A2(_01136_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06300_ (.A1(\as2650.instruction_args_latch[10] ),
    .A2(_01124_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06301_ (.A1(_01140_),
    .A2(_01144_),
    .A3(_01145_),
    .B(_01146_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06302_ (.A1(_00966_),
    .A2(_01127_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06303_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_01124_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06304_ (.A1(_01140_),
    .A2(_01148_),
    .B(_01149_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06305_ (.I(\as2650.instruction_args_latch[9] ),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06306_ (.I(_00967_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06307_ (.A1(_01128_),
    .A2(_01132_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06308_ (.A1(_01152_),
    .A2(_01134_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06309_ (.A1(_01151_),
    .A2(_01152_),
    .B1(_01153_),
    .B2(_01154_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06310_ (.A1(_01147_),
    .A2(_01150_),
    .A3(_01155_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06311_ (.A1(_01143_),
    .A2(_01156_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06312_ (.A1(_01113_),
    .A2(_01123_),
    .B(_01157_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06313_ (.I(_01129_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06314_ (.A1(\as2650.indirect_target[12] ),
    .A2(_01159_),
    .B1(_01137_),
    .B2(\as2650.PC[12] ),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06315_ (.A1(_01141_),
    .A2(_01160_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06316_ (.A1(\as2650.instruction_args_latch[12] ),
    .A2(_01140_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06317_ (.A1(_01125_),
    .A2(_01161_),
    .B(_01162_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06318_ (.A1(_01158_),
    .A2(_01163_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06319_ (.I(_00667_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06320_ (.I(_01165_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06321_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_01166_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06322_ (.A1(_00669_),
    .A2(_01164_),
    .B(_01167_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06323_ (.A1(\as2650.last_addr[12] ),
    .A2(_01168_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06324_ (.I(_00733_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06325_ (.A1(_01170_),
    .A2(_00731_),
    .B(_00748_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06326_ (.A1(_00733_),
    .A2(_00731_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06327_ (.A1(\as2650.page_reg[0] ),
    .A2(_01172_),
    .B(_01152_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06328_ (.A1(_01133_),
    .A2(_01135_),
    .A3(_01138_),
    .A4(_01160_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06329_ (.A1(\as2650.indirect_target[13] ),
    .A2(_01159_),
    .B1(_01137_),
    .B2(\as2650.page_reg[0] ),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06330_ (.A1(_01174_),
    .A2(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06331_ (.I(_01152_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06332_ (.A1(_01171_),
    .A2(_01173_),
    .B1(_01176_),
    .B2(_01177_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06333_ (.I(_01178_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06334_ (.A1(_01113_),
    .A2(_01123_),
    .B(_01157_),
    .C(_01163_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06335_ (.A1(_01179_),
    .A2(_01180_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06336_ (.A1(_00662_),
    .A2(_00676_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06337_ (.A1(_00659_),
    .A2(_01182_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06338_ (.I(_01183_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06339_ (.I(_01184_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06340_ (.A1(_01163_),
    .A2(_01178_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06341_ (.A1(_01112_),
    .A2(_01122_),
    .B(_01157_),
    .C(_01186_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06342_ (.A1(_01185_),
    .A2(_01187_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06343_ (.A1(\as2650.ivectors_base[9] ),
    .A2(_01166_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06344_ (.A1(_01181_),
    .A2(_01188_),
    .B(_01189_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06345_ (.A1(\as2650.last_addr[13] ),
    .A2(_01190_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06346_ (.A1(_01169_),
    .A2(_01191_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06347_ (.I(_01125_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06348_ (.A1(_01193_),
    .A2(_01144_),
    .A3(_01145_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06349_ (.A1(_01113_),
    .A2(_01123_),
    .B(_01150_),
    .C(_01155_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06350_ (.A1(_01146_),
    .A2(_01194_),
    .A3(_01195_),
    .Z(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06351_ (.I(_01183_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06352_ (.I(_01156_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06353_ (.A1(net308),
    .A2(_01123_),
    .B(_01198_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06354_ (.A1(_01197_),
    .A2(_01199_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06355_ (.A1(\as2650.ivectors_base[6] ),
    .A2(_00668_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06356_ (.A1(_01196_),
    .A2(_01200_),
    .B(_01201_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06357_ (.A1(\as2650.last_addr[10] ),
    .A2(_01202_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06358_ (.A1(_01199_),
    .A2(_01143_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06359_ (.I(_01165_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06360_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_01205_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06361_ (.A1(_00669_),
    .A2(_01204_),
    .B(_01206_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06362_ (.A1(_01207_),
    .A2(\as2650.last_addr[11] ),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _06363_ (.A1(_01113_),
    .A2(_01122_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06364_ (.A1(_01209_),
    .A2(_01150_),
    .B(_01155_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06365_ (.A1(_01197_),
    .A2(_01195_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06366_ (.A1(\as2650.ivectors_base[5] ),
    .A2(_01205_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06367_ (.A1(_01210_),
    .A2(_01211_),
    .B(_01212_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06368_ (.A1(\as2650.last_addr[9] ),
    .A2(_01213_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06369_ (.A1(_01209_),
    .A2(_01150_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06370_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_01166_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06371_ (.A1(_00669_),
    .A2(_01215_),
    .B(_01216_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06372_ (.A1(_01217_),
    .A2(\as2650.last_addr[8] ),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06373_ (.A1(_01203_),
    .A2(_01208_),
    .A3(_01214_),
    .A4(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06374_ (.I(_01166_),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06375_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_01220_),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06376_ (.I(_01172_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06377_ (.A1(\as2650.page_reg[1] ),
    .A2(_01172_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06378_ (.A1(_00756_),
    .A2(_01222_),
    .B(_01223_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06379_ (.I(_01175_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06380_ (.A1(_01174_),
    .A2(_01225_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06381_ (.I(_01137_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06382_ (.A1(\as2650.indirect_target[14] ),
    .A2(_01159_),
    .B1(_01227_),
    .B2(\as2650.page_reg[1] ),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06383_ (.A1(_01226_),
    .A2(_01228_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06384_ (.A1(_01226_),
    .A2(_01228_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06385_ (.A1(_01193_),
    .A2(_01230_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06386_ (.A1(_01193_),
    .A2(_01224_),
    .B1(_01229_),
    .B2(_01231_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06387_ (.I(_01177_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06388_ (.A1(\as2650.indirect_target[15] ),
    .A2(_01159_),
    .B1(_01227_),
    .B2(\as2650.page_reg[2] ),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06389_ (.A1(_01230_),
    .A2(_01234_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06390_ (.I0(\as2650.instruction_args_latch[15] ),
    .I1(\as2650.page_reg[2] ),
    .S(_01222_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06391_ (.A1(_01177_),
    .A2(_01236_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06392_ (.A1(_01233_),
    .A2(_01235_),
    .B(_01237_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06393_ (.A1(_01187_),
    .A2(_01232_),
    .A3(_01238_),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06394_ (.A1(_01187_),
    .A2(_01232_),
    .B(_01238_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06395_ (.A1(_01239_),
    .A2(_01240_),
    .B(_01220_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06396_ (.A1(_01221_),
    .A2(_01241_),
    .B(\as2650.last_addr[15] ),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06397_ (.A1(\as2650.last_addr[15] ),
    .A2(_01221_),
    .A3(_01241_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06398_ (.A1(_01187_),
    .A2(_01232_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06399_ (.A1(\as2650.ivectors_base[10] ),
    .A2(_00668_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06400_ (.A1(_01185_),
    .A2(_01244_),
    .B(_01245_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06401_ (.A1(\as2650.last_addr[14] ),
    .A2(_01246_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06402_ (.A1(_01242_),
    .A2(_01243_),
    .B(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06403_ (.A1(_01192_),
    .A2(_01219_),
    .A3(_01248_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06404_ (.I(_00683_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06405_ (.I(_00660_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06406_ (.A1(_01251_),
    .A2(_01182_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06407_ (.A1(_01250_),
    .A2(_00680_),
    .B(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06408_ (.A1(_01249_),
    .A2(_01253_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06409_ (.I(_01254_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06410_ (.I(_01255_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06411_ (.I(_01256_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06412_ (.I(_01257_),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06413_ (.A1(wb_reset_override),
    .A2(wb_reset_override_en),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06414_ (.A1(wb_reset_override_en),
    .A2(net33),
    .B(_01258_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06415_ (.A1(net58),
    .A2(_01259_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _06416_ (.I(_01260_),
    .ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06417_ (.I(_00755_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06418_ (.I(_01012_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06419_ (.A1(_01261_),
    .A2(_01262_),
    .A3(_01017_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06420_ (.I(_01035_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06421_ (.A1(_01261_),
    .A2(_01264_),
    .B(_01036_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06422_ (.A1(_01261_),
    .A2(_01264_),
    .A3(_01036_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06423_ (.A1(_01263_),
    .A2(_01265_),
    .B(_01266_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06424_ (.A1(_01067_),
    .A2(_01065_),
    .A3(_01267_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06425_ (.A1(\as2650.irqs_latch[6] ),
    .A2(\as2650.irqs_latch[7] ),
    .A3(_01184_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06426_ (.A1(\as2650.irqs_latch[4] ),
    .A2(\as2650.irqs_latch[5] ),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06427_ (.A1(\as2650.irqs_latch[2] ),
    .A2(\as2650.irqs_latch[3] ),
    .B(_01270_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06428_ (.A1(_01269_),
    .A2(_01271_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06429_ (.A1(_00668_),
    .A2(_01268_),
    .B(_01272_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06430_ (.A1(_01261_),
    .A2(_01262_),
    .B(_01017_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06431_ (.A1(_01018_),
    .A2(_01274_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06432_ (.A1(_00682_),
    .A2(_01183_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06433_ (.A1(_01184_),
    .A2(_01275_),
    .B(_01276_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06434_ (.A1(\as2650.last_addr[0] ),
    .A2(_01277_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06435_ (.A1(_01266_),
    .A2(_01034_),
    .B(_01018_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06436_ (.A1(_01037_),
    .A2(_01263_),
    .A3(_01265_),
    .B(_01183_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06437_ (.I(\as2650.irqs_latch[2] ),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06438_ (.A1(\as2650.irqs_latch[1] ),
    .A2(_01281_),
    .B(\as2650.irqs_latch[3] ),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06439_ (.A1(\as2650.irqs_latch[4] ),
    .A2(_01282_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06440_ (.A1(\as2650.irqs_latch[5] ),
    .A2(_01283_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06441_ (.A1(\as2650.irqs_latch[6] ),
    .A2(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06442_ (.A1(\as2650.irqs_latch[7] ),
    .A2(_01285_),
    .B(_00667_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06443_ (.A1(_01279_),
    .A2(_01280_),
    .B(_01286_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06444_ (.A1(\as2650.last_addr[1] ),
    .A2(_01287_),
    .Z(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06445_ (.A1(\as2650.last_addr[2] ),
    .A2(_01273_),
    .B(_01278_),
    .C(_01288_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06446_ (.A1(\as2650.last_addr[2] ),
    .A2(_01273_),
    .B(_01289_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06447_ (.A1(_01067_),
    .A2(_01065_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06448_ (.A1(_01067_),
    .A2(_01065_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06449_ (.A1(_01267_),
    .A2(_01291_),
    .B(_01292_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06450_ (.A1(_01293_),
    .A2(_01085_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06451_ (.A1(_01269_),
    .A2(_01270_),
    .B1(_01294_),
    .B2(_01197_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06452_ (.A1(\as2650.last_addr[3] ),
    .A2(_01295_),
    .Z(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06453_ (.A1(_01080_),
    .A2(_01084_),
    .Z(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06454_ (.A1(_01080_),
    .A2(_01084_),
    .Z(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06455_ (.A1(_01293_),
    .A2(_01297_),
    .B(_01298_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06456_ (.A1(_01299_),
    .A2(net314),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06457_ (.A1(_01299_),
    .A2(net314),
    .B(_01184_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06458_ (.A1(\as2650.ivectors_base[0] ),
    .A2(_01165_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06459_ (.A1(_01300_),
    .A2(_01301_),
    .B(_01302_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06460_ (.A1(\as2650.last_addr[4] ),
    .A2(_01303_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06461_ (.A1(_01290_),
    .A2(_01296_),
    .A3(_01304_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06462_ (.I(\as2650.ivectors_base[1] ),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06463_ (.A1(_01115_),
    .A2(_01300_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06464_ (.A1(_01101_),
    .A2(_01307_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06465_ (.I0(_01306_),
    .I1(_01308_),
    .S(_01197_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06466_ (.A1(\as2650.last_addr[5] ),
    .A2(_01309_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06467_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_01205_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06468_ (.A1(_00991_),
    .A2(_01118_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06469_ (.A1(_01087_),
    .A2(_01111_),
    .B(_01117_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06470_ (.A1(_01312_),
    .A2(_01313_),
    .B(_01165_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06471_ (.A1(_01312_),
    .A2(_01313_),
    .B(_01314_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06472_ (.A1(_01311_),
    .A2(_01315_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06473_ (.A1(\as2650.last_addr[6] ),
    .A2(_01316_),
    .Z(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06474_ (.A1(_01312_),
    .A2(_01313_),
    .B(_01119_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06475_ (.A1(_00974_),
    .A2(_01318_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06476_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_01205_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06477_ (.A1(_00669_),
    .A2(_01319_),
    .B(_01320_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06478_ (.A1(\as2650.last_addr[7] ),
    .A2(_01321_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06479_ (.A1(_01305_),
    .A2(_01310_),
    .A3(_01317_),
    .A4(_01322_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06480_ (.A1(_01253_),
    .A2(_01323_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06481_ (.A1(_01249_),
    .A2(_01324_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06482_ (.I(_01325_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06483_ (.I(_01326_),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06484_ (.I0(_01006_),
    .I1(_00999_),
    .S(_00582_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06485_ (.I(_01327_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06486_ (.I(_01328_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06487_ (.I(_01329_),
    .Z(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06488_ (.I(_01330_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06489_ (.I(_01331_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06490_ (.I(_01332_),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06491_ (.A1(_00581_),
    .A2(_00870_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06492_ (.A1(_00587_),
    .A2(_01025_),
    .B(_01333_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06493_ (.I(_01334_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06494_ (.I(_01335_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06495_ (.I(_01336_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06496_ (.I(_01337_),
    .Z(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06497_ (.I(_01338_),
    .Z(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06498_ (.I(_01339_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06499_ (.I(_01340_),
    .Z(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06500_ (.I(_01341_),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06501_ (.A1(_00581_),
    .A2(_00912_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06502_ (.A1(_00798_),
    .A2(_01046_),
    .B(_01342_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06503_ (.I(_01343_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06504_ (.I(_01344_),
    .Z(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06505_ (.I(_01345_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06506_ (.I(_01346_),
    .Z(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06507_ (.I(_01347_),
    .Z(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06508_ (.I(_01348_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06509_ (.I(_01349_),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06510_ (.I0(\as2650.regs[0][3] ),
    .I1(\as2650.regs[4][3] ),
    .S(_00620_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06511_ (.I(_01350_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06512_ (.I(_01351_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06513_ (.I(_01352_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06514_ (.I(_01353_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06515_ (.I(_01354_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06516_ (.I(_01355_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06517_ (.I(_01356_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06518_ (.I(_01357_),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _06519_ (.I(wb_io3_test),
    .ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06520_ (.A1(_01192_),
    .A2(_01219_),
    .A3(_01248_),
    .A4(_01323_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06521_ (.I(_01358_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06522_ (.I(_01359_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06523_ (.I(_01360_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06524_ (.I(_01361_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _06525_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net215),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06526_ (.I(_01363_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06527_ (.I(_01364_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06528_ (.I(_01365_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06529_ (.I(_01366_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06530_ (.I(_01367_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06531_ (.I(_00682_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06532_ (.I(_01369_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06533_ (.A1(_00722_),
    .A2(_00726_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06534_ (.I(_01371_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06535_ (.I(_01372_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06536_ (.I(_01373_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06537_ (.I(_00659_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06538_ (.A1(_01375_),
    .A2(_00666_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06539_ (.A1(_00716_),
    .A2(_00719_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06540_ (.I(_01377_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06541_ (.I(_01378_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06542_ (.A1(_00735_),
    .A2(_00736_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06543_ (.I(_00721_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06544_ (.I(_00711_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06545_ (.A1(net40),
    .A2(_01382_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06546_ (.A1(net52),
    .A2(_00743_),
    .B(_01383_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06547_ (.A1(\as2650.insin[2] ),
    .A2(_00721_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06548_ (.A1(_01381_),
    .A2(_01384_),
    .B(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06549_ (.A1(_01380_),
    .A2(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06550_ (.I(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06551_ (.I(_01388_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06552_ (.I(_01389_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06553_ (.I(_01390_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06554_ (.I(_01391_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06555_ (.I(_01392_),
    .Z(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06556_ (.I(_00731_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06557_ (.A1(_00709_),
    .A2(_00715_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06558_ (.I(_01395_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06559_ (.A1(_01394_),
    .A2(_01396_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06560_ (.A1(_01393_),
    .A2(_01397_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06561_ (.A1(_01379_),
    .A2(_01398_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06562_ (.A1(_01376_),
    .A2(_01399_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06563_ (.A1(_01374_),
    .A2(_01400_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06564_ (.I(_00675_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06565_ (.I(_00662_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06566_ (.A1(_01369_),
    .A2(_01403_),
    .A3(_00941_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06567_ (.I(_01404_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06568_ (.A1(_01402_),
    .A2(_01405_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06569_ (.A1(_00700_),
    .A2(_00707_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06570_ (.A1(_01371_),
    .A2(_01407_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06571_ (.A1(_00745_),
    .A2(_00746_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06572_ (.A1(_00716_),
    .A2(_00719_),
    .Z(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06573_ (.I(_01410_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06574_ (.A1(_01409_),
    .A2(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06575_ (.I(_00892_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06576_ (.I(_01413_),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06577_ (.I(_01414_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06578_ (.I(_01415_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06579_ (.A1(_00695_),
    .A2(_00698_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06580_ (.A1(_00728_),
    .A2(_00729_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06581_ (.A1(_01417_),
    .A2(_01418_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06582_ (.A1(_01394_),
    .A2(_01419_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06583_ (.A1(_01412_),
    .A2(_01416_),
    .A3(_01392_),
    .A4(_01420_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06584_ (.I(_01394_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06585_ (.I(_00737_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06586_ (.I(_01423_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06587_ (.I(_01409_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06588_ (.A1(_01422_),
    .A2(_01424_),
    .B(_01425_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06589_ (.A1(_01379_),
    .A2(_01408_),
    .A3(_01421_),
    .A4(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06590_ (.I(_01427_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06591_ (.I(_01428_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06592_ (.A1(_01233_),
    .A2(_01406_),
    .B(_01429_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06593_ (.A1(_01370_),
    .A2(_01401_),
    .B(_01430_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06594_ (.A1(_01252_),
    .A2(_01362_),
    .B(_01368_),
    .C(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06595_ (.I(net260),
    .ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06596_ (.I(_01382_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06597_ (.I(_01433_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06598_ (.I(_01434_),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06599_ (.I(\as2650.io_bus_we ),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06600_ (.I(\as2650.ext_io_addr[7] ),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06601_ (.I(_01436_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06602_ (.I(\as2650.ext_io_addr[6] ),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06603_ (.I(_01438_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06604_ (.A1(_01435_),
    .A2(_01437_),
    .A3(_01439_),
    .ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06605_ (.I(_01437_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06606_ (.A1(\as2650.io_bus_we ),
    .A2(_01440_),
    .A3(_01439_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06607_ (.I(_01441_),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06608_ (.A1(_01435_),
    .A2(_01440_),
    .A3(_01439_),
    .ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06609_ (.A1(\as2650.io_bus_we ),
    .A2(_01437_),
    .A3(_01439_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06610_ (.I(_01442_),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06611_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .A3(net215),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06612_ (.I(_01443_),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06613_ (.I(_01444_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06614_ (.I(_01445_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06615_ (.I(_01446_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06616_ (.I(_01447_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06617_ (.I(_01448_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06618_ (.I(_01449_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06619_ (.I(_01256_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06620_ (.I(_01401_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06621_ (.A1(_01451_),
    .A2(_01326_),
    .A3(_01452_),
    .A4(net260),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06622_ (.A1(_01450_),
    .A2(_01453_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06623_ (.A1(_01250_),
    .A2(_00680_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06624_ (.I(_01362_),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06625_ (.I(_01417_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06626_ (.I(_01456_),
    .Z(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06627_ (.I(_01457_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _06628_ (.A1(_01454_),
    .A2(_01455_),
    .B1(_01400_),
    .B2(_01458_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06629_ (.I(_01368_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06630_ (.A1(_01460_),
    .A2(_01430_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06631_ (.A1(_01459_),
    .A2(_01461_),
    .ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06632_ (.I(_01447_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06633_ (.I(_01462_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06634_ (.A1(clknet_leaf_59_wb_clk_i),
    .A2(net213),
    .A3(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06635_ (.I(_01464_),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06636_ (.A1(clknet_leaf_59_wb_clk_i),
    .A2(net214),
    .A3(_01463_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06637_ (.I(_01465_),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06638_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_159_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06639_ (.A1(\web_behavior[1] ),
    .A2(clknet_leaf_159_wb_clk_i),
    .B(\web_behavior[0] ),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06640__1 (.I(_01467_),
    .ZN(net303));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06641_ (.A1(_01466_),
    .A2(net303),
    .B(_01432_),
    .ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06642_ (.I(wb_debug_carry),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _06643_ (.I(\as2650.debug_psl[0] ),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06644_ (.I(\as2650.debug_psl[6] ),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06645_ (.I(_01471_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06646_ (.I(_01472_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06647_ (.I(_01418_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06648_ (.I(_01474_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06649_ (.I(_01475_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06650_ (.A1(wb_debug_cc),
    .A2(_01252_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06651_ (.A1(wb_debug_cc),
    .A2(_01473_),
    .B1(_01476_),
    .B2(_01477_),
    .C(wb_debug_carry),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06652_ (.A1(_01469_),
    .A2(_01470_),
    .B(_01478_),
    .ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06653_ (.I(\as2650.debug_psl[7] ),
    .Z(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06654_ (.I(_01479_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06655_ (.I(_01407_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06656_ (.A1(wb_debug_cc),
    .A2(_01480_),
    .B1(_01481_),
    .B2(_01477_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06657_ (.I(\as2650.debug_psl[5] ),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06658_ (.I(_01483_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06659_ (.I(_01484_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06660_ (.I(_01485_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06661_ (.A1(_01469_),
    .A2(_01486_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06662_ (.A1(_01469_),
    .A2(_01482_),
    .B(_01487_),
    .ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06663_ (.I(_00597_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06664_ (.I(_01488_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06665_ (.I(_01489_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06666_ (.I(_01490_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06667_ (.I(_01491_),
    .Z(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06668_ (.I(_01492_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06669_ (.I(_01493_),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06670_ (.I(_01494_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06671_ (.I(_01493_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06672_ (.A1(_01496_),
    .A2(\as2650.regs[6][0] ),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06673_ (.A1(_01495_),
    .A2(_00885_),
    .B(_01497_),
    .ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06674_ (.A1(_01496_),
    .A2(\as2650.regs[6][1] ),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06675_ (.A1(_01495_),
    .A2(_00872_),
    .B(_01498_),
    .ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06676_ (.I(_01493_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06677_ (.A1(_01499_),
    .A2(\as2650.regs[6][2] ),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06678_ (.A1(_01495_),
    .A2(_00914_),
    .B(_01500_),
    .ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06679_ (.A1(_01499_),
    .A2(\as2650.regs[6][3] ),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06680_ (.A1(_01495_),
    .A2(_00902_),
    .B(_01501_),
    .ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06681_ (.A1(_01499_),
    .A2(\as2650.regs[6][4] ),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06682_ (.A1(_01496_),
    .A2(_00852_),
    .B(_01502_),
    .ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06683_ (.A1(_01499_),
    .A2(\as2650.regs[6][5] ),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06684_ (.A1(_01496_),
    .A2(_00836_),
    .B(_01503_),
    .ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06685_ (.I0(\as2650.regs[2][6] ),
    .I1(\as2650.regs[6][6] ),
    .S(_01494_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06686_ (.I(_01504_),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06687_ (.I0(\as2650.regs[2][7] ),
    .I1(\as2650.regs[6][7] ),
    .S(_01494_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06688_ (.I(_01505_),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06689_ (.I(_00597_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06690_ (.A1(_01506_),
    .A2(\as2650.regs[7][0] ),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06691_ (.A1(_01488_),
    .A2(_01002_),
    .B(_01507_),
    .ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06692_ (.A1(_01506_),
    .A2(\as2650.regs[7][1] ),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06693_ (.A1(_01488_),
    .A2(_01022_),
    .B(_01508_),
    .ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06694_ (.A1(_01488_),
    .A2(\as2650.regs[7][2] ),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06695_ (.A1(_01489_),
    .A2(_01043_),
    .B(_01509_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06696_ (.I(_01510_),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06697_ (.I0(\as2650.regs[3][3] ),
    .I1(\as2650.regs[7][3] ),
    .S(_01506_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06698_ (.I(_01511_),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06699_ (.I(_00626_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06700_ (.I(_01512_),
    .Z(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06701_ (.A1(_01512_),
    .A2(\as2650.regs[3][4] ),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06702_ (.A1(_01513_),
    .A2(_00844_),
    .B(_01514_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06703_ (.I(_01515_),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06704_ (.A1(_01512_),
    .A2(\as2650.regs[3][5] ),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06705_ (.A1(_01512_),
    .A2(_00827_),
    .B(_01516_),
    .ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06706_ (.I0(\as2650.regs[3][6] ),
    .I1(\as2650.regs[7][6] ),
    .S(_01489_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _06707_ (.I(_01517_),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06708_ (.I0(\as2650.regs[3][7] ),
    .I1(\as2650.regs[7][7] ),
    .S(_01489_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06709_ (.I(_01518_),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06710_ (.I(_01422_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06711_ (.A1(_00789_),
    .A2(_01001_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06712_ (.I(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06713_ (.I(_01521_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06714_ (.A1(_01395_),
    .A2(_01410_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06715_ (.A1(_01391_),
    .A2(_01523_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06716_ (.A1(_01456_),
    .A2(_01474_),
    .A3(_01524_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06717_ (.I(_01525_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06718_ (.A1(_01519_),
    .A2(_01522_),
    .A3(_01526_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06719_ (.I(_01527_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06720_ (.A1(_01359_),
    .A2(_01381_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06721_ (.A1(_01528_),
    .A2(_01529_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06722_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06723_ (.A1(_01366_),
    .A2(_01531_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06724_ (.I(_01532_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06725_ (.I(_01529_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06726_ (.A1(\as2650.chirp_ptr[1] ),
    .A2(\as2650.chirp_ptr[0] ),
    .A3(_01528_),
    .A4(_01533_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06727_ (.A1(\as2650.chirp_ptr[2] ),
    .A2(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06728_ (.I(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06729_ (.A1(_01447_),
    .A2(_01535_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06730_ (.I(_01537_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06731_ (.I(_01538_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06732_ (.I(_00373_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06733_ (.A1(\as2650.chirp_ptr[0] ),
    .A2(_01528_),
    .A3(_01533_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06734_ (.A1(\as2650.chirp_ptr[1] ),
    .A2(_01540_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06735_ (.A1(_01447_),
    .A2(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06736_ (.A1(_01539_),
    .A2(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06737_ (.A1(_01531_),
    .A2(_01542_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06738_ (.A1(_01543_),
    .A2(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06739_ (.A1(_00373_),
    .A2(_01536_),
    .B1(_00375_),
    .B2(_01545_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06740_ (.A1(_01539_),
    .A2(_01537_),
    .A3(_01542_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06741_ (.A1(_01544_),
    .A2(_01546_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06742_ (.A1(_01538_),
    .A2(_01541_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06743_ (.A1(_00375_),
    .A2(_01545_),
    .B(_01547_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06744_ (.A1(_01537_),
    .A2(_01544_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(_01538_),
    .A2(_01543_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06746_ (.A1(_01548_),
    .A2(_00116_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06747_ (.I(_01549_),
    .Z(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06748_ (.A1(_01546_),
    .A2(_01547_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06749_ (.I(_01550_),
    .Z(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06750_ (.I(_01325_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06751_ (.I(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06752_ (.A1(_00685_),
    .A2(_00752_),
    .B(_01177_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06753_ (.A1(_01009_),
    .A2(_01553_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06754_ (.I(_00685_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06755_ (.A1(_00732_),
    .A2(_00742_),
    .A3(_00751_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06756_ (.A1(_01555_),
    .A2(_01556_),
    .B(_01125_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06757_ (.I(_01329_),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06758_ (.A1(_00892_),
    .A2(_01558_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06759_ (.A1(_00892_),
    .A2(_01262_),
    .B(_01557_),
    .C(_01559_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06760_ (.A1(_01554_),
    .A2(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06761_ (.A1(_01217_),
    .A2(_01257_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06762_ (.A1(_01451_),
    .A2(_01561_),
    .B(_01562_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06763_ (.A1(_01552_),
    .A2(_01563_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06764_ (.I(_01326_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06765_ (.A1(_01277_),
    .A2(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06766_ (.A1(_01564_),
    .A2(_01566_),
    .ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06767_ (.I(_01051_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06768_ (.I(_01567_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06769_ (.I(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06770_ (.I(_01452_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06771_ (.I(_01325_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06772_ (.I(_01256_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06773_ (.I(_01553_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06774_ (.A1(_01051_),
    .A2(_01573_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06775_ (.I(_01557_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06776_ (.A1(_01413_),
    .A2(_01339_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06777_ (.A1(_01414_),
    .A2(net309),
    .B(_01575_),
    .C(_01576_),
    .ZN(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06778_ (.A1(_01574_),
    .A2(_01577_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06779_ (.I(_01255_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06780_ (.A1(_01213_),
    .A2(_01579_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06781_ (.A1(_01572_),
    .A2(_01578_),
    .B(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06782_ (.A1(_01571_),
    .A2(_01581_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06783_ (.I(_01326_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06784_ (.I(_01401_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06785_ (.A1(_01287_),
    .A2(_01583_),
    .B(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06786_ (.A1(_01569_),
    .A2(_01570_),
    .B1(_01582_),
    .B2(_01585_),
    .ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06787_ (.I(_01053_),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06788_ (.I(_01586_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06789_ (.I(_01587_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06790_ (.I(_01325_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06791_ (.I(_00989_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06792_ (.A1(_01590_),
    .A2(_01056_),
    .A3(_01058_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06793_ (.A1(_01590_),
    .A2(_01055_),
    .B(_01591_),
    .C(_01413_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06794_ (.I(_00797_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06795_ (.I(_01343_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06796_ (.A1(_01593_),
    .A2(_01594_),
    .B(_01557_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06797_ (.A1(_01048_),
    .A2(_01575_),
    .B1(_01592_),
    .B2(_01595_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(_01202_),
    .A2(_01256_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06799_ (.A1(_01257_),
    .A2(_01596_),
    .B(_01597_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06800_ (.A1(_01273_),
    .A2(_01551_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06801_ (.A1(_01589_),
    .A2(_01598_),
    .B(_01599_),
    .C(_01452_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06802_ (.A1(_01588_),
    .A2(_01570_),
    .B(_01600_),
    .ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06803_ (.I(_01070_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06804_ (.I(_01601_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06805_ (.I(_01602_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06806_ (.A1(_01413_),
    .A2(_01354_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06807_ (.A1(_01593_),
    .A2(_01074_),
    .A3(_01079_),
    .B(_01604_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06808_ (.I0(_01070_),
    .I1(_01605_),
    .S(_01553_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06809_ (.A1(_01207_),
    .A2(_01579_),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06810_ (.A1(_01572_),
    .A2(_01606_),
    .B(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06811_ (.A1(_01571_),
    .A2(_01608_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06812_ (.A1(_01295_),
    .A2(_01583_),
    .B(_01584_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06813_ (.A1(_01603_),
    .A2(_01570_),
    .B1(_01609_),
    .B2(_01610_),
    .ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06814_ (.I(_01093_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06815_ (.I(_01611_),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06816_ (.I(_01612_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06817_ (.A1(_01039_),
    .A2(_01104_),
    .B(_01106_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06818_ (.I(_00653_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06819_ (.A1(_01615_),
    .A2(_01414_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06820_ (.A1(_01414_),
    .A2(_01614_),
    .B(_01616_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06821_ (.I0(_01093_),
    .I1(_01617_),
    .S(_01573_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06822_ (.I(_01618_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06823_ (.A1(_01168_),
    .A2(_01579_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06824_ (.A1(_01572_),
    .A2(_01619_),
    .B(_01620_),
    .ZN(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06825_ (.A1(_01589_),
    .A2(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06826_ (.A1(_01303_),
    .A2(_01565_),
    .B(_01584_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06827_ (.A1(_01613_),
    .A2(_01570_),
    .B1(_01622_),
    .B2(_01623_),
    .ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06828_ (.A1(_00833_),
    .A2(_00835_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06829_ (.A1(_00838_),
    .A2(_00841_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06830_ (.A1(_01624_),
    .A2(_01625_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06831_ (.I(_01575_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06832_ (.I(_01627_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06833_ (.A1(_00987_),
    .A2(_01094_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06834_ (.I0(_01092_),
    .I1(_01629_),
    .S(_01590_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06835_ (.A1(_01415_),
    .A2(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06836_ (.I(_00645_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06837_ (.I(_01593_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06838_ (.A1(_01632_),
    .A2(_01633_),
    .B(_01627_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06839_ (.A1(_01626_),
    .A2(_01628_),
    .B1(_01631_),
    .B2(_01634_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06840_ (.I(_01635_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06841_ (.A1(_01190_),
    .A2(_01257_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06842_ (.A1(_01451_),
    .A2(_01636_),
    .B(_01637_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06843_ (.A1(_01552_),
    .A2(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06844_ (.A1(_01309_),
    .A2(_01551_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06845_ (.A1(_01639_),
    .A2(_01640_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06846_ (.I(_00984_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06847_ (.I(_01641_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06848_ (.I(_01254_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06849_ (.A1(_01246_),
    .A2(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06850_ (.A1(_00641_),
    .A2(_01415_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06851_ (.A1(_01415_),
    .A2(_00990_),
    .B(_01627_),
    .C(_01645_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06852_ (.A1(_00929_),
    .A2(_01628_),
    .B(_01646_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06853_ (.I(_01647_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06854_ (.A1(_01572_),
    .A2(_01648_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06855_ (.A1(_01644_),
    .A2(_01649_),
    .B(_01589_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06856_ (.A1(_01316_),
    .A2(_01565_),
    .B(_01452_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06857_ (.A1(_01642_),
    .A2(_01584_),
    .B1(_01650_),
    .B2(_01651_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06858_ (.I(_01628_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06859_ (.I(_00628_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06860_ (.A1(_00924_),
    .A2(_00936_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06861_ (.A1(_01633_),
    .A2(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06862_ (.A1(_01653_),
    .A2(_01633_),
    .B(_01628_),
    .C(_01655_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06863_ (.A1(_00808_),
    .A2(_01652_),
    .B(_01656_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06864_ (.I(_01657_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06865_ (.A1(_01221_),
    .A2(_01241_),
    .B(_01579_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06866_ (.A1(_01451_),
    .A2(_01658_),
    .B(_01659_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06867_ (.A1(_01552_),
    .A2(_01660_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06868_ (.A1(_01321_),
    .A2(_01565_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06869_ (.A1(_01661_),
    .A2(_01662_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _06870_ (.A1(_01192_),
    .A2(_01219_),
    .A3(_01248_),
    .A4(_01323_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06871_ (.I(_01663_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06872_ (.I(_01664_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06873_ (.A1(_01665_),
    .A2(_01405_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06874_ (.A1(_01394_),
    .A2(_01386_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06875_ (.I(_01667_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06876_ (.A1(_01424_),
    .A2(_01668_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06877_ (.A1(_01170_),
    .A2(_01669_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06878_ (.I(_00741_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06879_ (.A1(_01380_),
    .A2(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06880_ (.A1(_01402_),
    .A2(_01672_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06881_ (.A1(_01670_),
    .A2(_01673_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06882_ (.A1(_01666_),
    .A2(_01674_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06883_ (.I(_01675_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06884_ (.A1(net36),
    .A2(_00743_),
    .B(_00691_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06885_ (.I(_01677_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06886_ (.A1(_01663_),
    .A2(_01443_),
    .A3(_01404_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06887_ (.I(_01679_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06888_ (.A1(\as2650.instruction_args_latch[15] ),
    .A2(_01679_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06889_ (.A1(_01678_),
    .A2(_01680_),
    .B(_01681_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06890_ (.A1(_01222_),
    .A2(_01682_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06891_ (.A1(_01424_),
    .A2(_01386_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06892_ (.A1(_01684_),
    .A2(_01683_),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06893_ (.A1(_01425_),
    .A2(_01685_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06894_ (.A1(_01676_),
    .A2(_01686_),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06895_ (.I(_01666_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06896_ (.I(_01688_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06897_ (.A1(_01402_),
    .A2(_01381_),
    .A3(_01689_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06898_ (.I(_01368_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06899_ (.I(_01691_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06900_ (.A1(_01687_),
    .A2(_01690_),
    .B(_01692_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06901_ (.I(net58),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06902_ (.I(net62),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06903_ (.I(net61),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06904_ (.A1(_01693_),
    .A2(_01694_),
    .A3(_01695_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06905_ (.A1(net96),
    .A2(net63),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06906_ (.A1(wb_feedback_delay),
    .A2(_01697_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06907_ (.A1(net97),
    .A2(_01698_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06908_ (.I(net59),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06909_ (.A1(_01700_),
    .A2(net60),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06910_ (.A1(_01699_),
    .A2(_01701_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06911_ (.A1(_01696_),
    .A2(net383),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06912_ (.I(net384),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06913_ (.I(_01704_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06914_ (.I0(net64),
    .I1(net114),
    .S(_01705_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06915_ (.I(_01706_),
    .Z(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06916_ (.I0(net75),
    .I1(net121),
    .S(_01705_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06917_ (.I(_01707_),
    .Z(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06918_ (.I0(net86),
    .I1(net122),
    .S(_01705_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06919_ (.I(_01708_),
    .Z(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06920_ (.I0(net89),
    .I1(net123),
    .S(_01705_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06921_ (.I(_01709_),
    .Z(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06922_ (.I(_01704_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06923_ (.I0(net90),
    .I1(net124),
    .S(_01710_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06924_ (.I(_01711_),
    .Z(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06925_ (.I0(net91),
    .I1(net125),
    .S(_01710_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06926_ (.I(_01712_),
    .Z(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06927_ (.I0(net92),
    .I1(net126),
    .S(_01710_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06928_ (.I(_01713_),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06929_ (.I0(net93),
    .I1(net127),
    .S(_01710_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06930_ (.I(_01714_),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06931_ (.I(_01704_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06932_ (.I0(net94),
    .I1(net128),
    .S(_01715_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06933_ (.I(_01716_),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06934_ (.I0(net95),
    .I1(net129),
    .S(_01715_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06935_ (.I(_01717_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06936_ (.I0(net65),
    .I1(net115),
    .S(_01715_),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06937_ (.I(_01718_),
    .Z(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06938_ (.I0(net66),
    .I1(net116),
    .S(_01715_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06939_ (.I(_01719_),
    .Z(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06940_ (.I(_01704_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06941_ (.I0(net67),
    .I1(net117),
    .S(_01720_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06942_ (.I(_01721_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06943_ (.I0(net68),
    .I1(net118),
    .S(_01720_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06944_ (.I(_01722_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06945_ (.I0(net69),
    .I1(net119),
    .S(_01720_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06946_ (.I(_01723_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06947_ (.I0(net70),
    .I1(net120),
    .S(_01720_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06948_ (.I(net385),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06949_ (.I(_01703_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06950_ (.I(_01725_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06951_ (.I0(net374),
    .I1(net98),
    .S(_01726_),
    .Z(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06952_ (.I(net375),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06953_ (.I0(net72),
    .I1(net105),
    .S(_01726_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06954_ (.I(_01728_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06955_ (.I0(net73),
    .I1(net106),
    .S(_01726_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06956_ (.I(_01729_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06957_ (.I0(net74),
    .I1(net107),
    .S(_01726_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06958_ (.I(_01730_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06959_ (.I(_01725_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06960_ (.I0(net76),
    .I1(net108),
    .S(_01731_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06961_ (.I(_01732_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06962_ (.I0(net77),
    .I1(net109),
    .S(_01731_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06963_ (.I(_01733_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06964_ (.I0(net78),
    .I1(net110),
    .S(_01731_),
    .Z(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06965_ (.I(_01734_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06966_ (.I0(net79),
    .I1(net111),
    .S(_01731_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06967_ (.I(_01735_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06968_ (.I(_01725_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06969_ (.I0(net80),
    .I1(net112),
    .S(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06970_ (.I(_01737_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06971_ (.I0(net81),
    .I1(net113),
    .S(_01736_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06972_ (.I(_01738_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06973_ (.I0(net82),
    .I1(net99),
    .S(_01736_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06974_ (.I(_01739_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06975_ (.I0(net83),
    .I1(net100),
    .S(_01736_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06976_ (.I(_01740_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06977_ (.I(_01725_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06978_ (.I0(net84),
    .I1(net101),
    .S(_01741_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06979_ (.I(_01742_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06980_ (.I0(net85),
    .I1(net102),
    .S(_01741_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06981_ (.I(_01743_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06982_ (.I0(net87),
    .I1(net103),
    .S(_01741_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06983_ (.I(_01744_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06984_ (.I0(net88),
    .I1(net104),
    .S(_01741_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06985_ (.I(_01745_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06986_ (.I(_01693_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06987_ (.I(net62),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06988_ (.I(_01747_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06989_ (.I(net59),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06990_ (.I(net60),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06991_ (.I(_01695_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06992_ (.A1(_01694_),
    .A2(_01699_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06993_ (.A1(_01749_),
    .A2(_01750_),
    .A3(_01751_),
    .A4(_01752_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06994_ (.A1(_01746_),
    .A2(_01748_),
    .A3(net401),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06995_ (.I0(net151),
    .I1(net64),
    .S(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06996_ (.I(_01755_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06997_ (.I0(net152),
    .I1(net75),
    .S(_01754_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06998_ (.I(_01756_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06999_ (.I0(net153),
    .I1(net86),
    .S(_01754_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07000_ (.I(_01757_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07001_ (.I(_01693_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07002_ (.I(_01758_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07003_ (.I(_01759_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07004_ (.A1(_01760_),
    .A2(wb_feedback_delay),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07005_ (.I(_01761_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07006_ (.A1(wb_feedback_delay),
    .A2(_01697_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07007_ (.I(_01762_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07008_ (.I(_01763_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07009_ (.A1(net225),
    .A2(_01764_),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07010_ (.I(_01747_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07011_ (.I(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07012_ (.I(net61),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07013_ (.I(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07014_ (.A1(_01700_),
    .A2(net114),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07015_ (.A1(_01750_),
    .A2(_01751_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07016_ (.A1(_01749_),
    .A2(net151),
    .B(_01771_),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07017_ (.A1(_01769_),
    .A2(_01470_),
    .B1(_01770_),
    .B2(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07018_ (.I(_01748_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07019_ (.I(\wb_counter[0] ),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07020_ (.A1(_01774_),
    .A2(_01775_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07021_ (.I(_01698_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07022_ (.A1(_01767_),
    .A2(_01773_),
    .B(_01776_),
    .C(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07023_ (.I(_01746_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07024_ (.I(_01779_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07025_ (.A1(_01765_),
    .A2(_01778_),
    .B(_01780_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07026_ (.A1(net236),
    .A2(_01764_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _07027_ (.I(\as2650.debug_psl[1] ),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07028_ (.A1(_01700_),
    .A2(net121),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07029_ (.A1(_01749_),
    .A2(net152),
    .B(_01771_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07030_ (.A1(_01769_),
    .A2(_01782_),
    .B1(_01783_),
    .B2(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07031_ (.I(_01694_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07032_ (.I(_01786_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07033_ (.I(\wb_counter[1] ),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07034_ (.A1(_01787_),
    .A2(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07035_ (.A1(_01767_),
    .A2(_01785_),
    .B(_01789_),
    .C(_01777_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07036_ (.A1(_01781_),
    .A2(_01790_),
    .B(_01780_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07037_ (.A1(net247),
    .A2(_01764_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07038_ (.I(\as2650.debug_psl[2] ),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07039_ (.I(_01792_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07040_ (.A1(_01700_),
    .A2(net122),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07041_ (.A1(_01749_),
    .A2(net153),
    .B(_01771_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07042_ (.A1(_01769_),
    .A2(_01793_),
    .B1(_01794_),
    .B2(_01795_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07043_ (.I(\wb_counter[2] ),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07044_ (.A1(_01787_),
    .A2(_01797_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07045_ (.A1(_01767_),
    .A2(_01796_),
    .B(_01798_),
    .C(_01777_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07046_ (.A1(_01791_),
    .A2(_01799_),
    .B(_01780_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07047_ (.I(_01693_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07048_ (.I(_01800_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07049_ (.I(_01762_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07050_ (.I(_01802_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07051_ (.I(\wb_counter[3] ),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07052_ (.I(net382),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07053_ (.I(_01805_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07054_ (.A1(net59),
    .A2(_01750_),
    .B(_01695_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07055_ (.I(_01807_),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07056_ (.A1(net123),
    .A2(_01806_),
    .B(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07057_ (.I(\as2650.debug_psl[3] ),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07058_ (.I(_01810_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07059_ (.I(_01811_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07060_ (.I(_01747_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07061_ (.A1(_01769_),
    .A2(_01812_),
    .B(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07062_ (.I(_01762_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07063_ (.I(_01815_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07064_ (.A1(_01787_),
    .A2(_01804_),
    .B1(_01809_),
    .B2(_01814_),
    .C(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07065_ (.A1(net250),
    .A2(_01803_),
    .B(_01817_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07066_ (.A1(_01801_),
    .A2(_01818_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07067_ (.I(\wb_counter[4] ),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07068_ (.A1(net124),
    .A2(_01806_),
    .B(_01808_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07069_ (.I(_01695_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07070_ (.I(_01786_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07071_ (.A1(_01492_),
    .A2(_01821_),
    .B(_01822_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07072_ (.A1(_01787_),
    .A2(_01819_),
    .B1(_01820_),
    .B2(_01823_),
    .C(_01816_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07073_ (.A1(net251),
    .A2(_01803_),
    .B(_01824_),
    .ZN(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07074_ (.A1(_01801_),
    .A2(_01825_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07075_ (.I(_01746_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07076_ (.I(_01826_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07077_ (.I(_01748_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07078_ (.I(\wb_counter[5] ),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07079_ (.A1(net125),
    .A2(_01806_),
    .B(_01808_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07080_ (.I(_01768_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07081_ (.A1(_01831_),
    .A2(_01486_),
    .B(_01822_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07082_ (.A1(_01828_),
    .A2(_01829_),
    .B1(_01830_),
    .B2(_01832_),
    .C(_01816_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07083_ (.A1(net252),
    .A2(_01803_),
    .B(_01833_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07084_ (.A1(_01827_),
    .A2(_01834_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07085_ (.I(\wb_counter[6] ),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07086_ (.A1(net126),
    .A2(_01806_),
    .B(_01808_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07087_ (.A1(_01473_),
    .A2(_01821_),
    .B(_01822_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07088_ (.A1(_01828_),
    .A2(_01835_),
    .B1(_01836_),
    .B2(_01837_),
    .C(_01816_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07089_ (.A1(net253),
    .A2(_01803_),
    .B(_01838_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07090_ (.A1(_01827_),
    .A2(_01839_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07091_ (.I(_01802_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07092_ (.I(\wb_counter[7] ),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07093_ (.I(_01805_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07094_ (.I(_01807_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07095_ (.A1(net127),
    .A2(_01842_),
    .B(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07096_ (.A1(_01480_),
    .A2(_01821_),
    .B(_01822_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07097_ (.I(_01815_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07098_ (.A1(_01828_),
    .A2(_01841_),
    .B1(_01844_),
    .B2(_01845_),
    .C(_01846_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07099_ (.A1(net254),
    .A2(_01840_),
    .B(_01847_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07100_ (.A1(_01827_),
    .A2(_01848_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07101_ (.I(\wb_counter[8] ),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07102_ (.A1(net128),
    .A2(_01842_),
    .B(_01843_),
    .ZN(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07103_ (.I(\as2650.debug_psu[0] ),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07104_ (.I(_01851_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07105_ (.I(_01786_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07106_ (.A1(_01831_),
    .A2(_01852_),
    .B(_01853_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07107_ (.A1(_01828_),
    .A2(_01849_),
    .B1(_01850_),
    .B2(_01854_),
    .C(_01846_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07108_ (.A1(net255),
    .A2(_01840_),
    .B(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07109_ (.A1(_01827_),
    .A2(_01856_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07110_ (.I(_01779_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07111_ (.I(_01748_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07112_ (.I(\wb_counter[9] ),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07113_ (.A1(net129),
    .A2(_01842_),
    .B(_01843_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07114_ (.I(\as2650.debug_psu[1] ),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07115_ (.I(_01861_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07116_ (.A1(_01831_),
    .A2(_01862_),
    .B(_01853_),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07117_ (.A1(_01858_),
    .A2(_01859_),
    .B1(_01860_),
    .B2(_01863_),
    .C(_01846_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07118_ (.A1(net256),
    .A2(_01840_),
    .B(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07119_ (.A1(_01857_),
    .A2(_01865_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07120_ (.I(\wb_counter[10] ),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07121_ (.A1(net115),
    .A2(_01842_),
    .B(_01843_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07122_ (.I(\as2650.debug_psu[2] ),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07123_ (.I(_01868_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07124_ (.I(_01869_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07125_ (.I(_01870_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07126_ (.A1(_01831_),
    .A2(_01871_),
    .B(_01853_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07127_ (.A1(_01858_),
    .A2(_01866_),
    .B1(_01867_),
    .B2(_01872_),
    .C(_01846_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07128_ (.A1(net226),
    .A2(_01840_),
    .B(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07129_ (.A1(_01857_),
    .A2(_01874_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07130_ (.I(_01802_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07131_ (.I(\wb_counter[11] ),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07132_ (.I(_01805_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07133_ (.I(_01807_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07134_ (.A1(net116),
    .A2(_01877_),
    .B(_01878_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07135_ (.I(_01768_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07136_ (.I(\as2650.debug_psu[3] ),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07137_ (.I(_01881_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07138_ (.A1(_01880_),
    .A2(_01882_),
    .B(_01853_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07139_ (.I(_01762_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07140_ (.A1(_01858_),
    .A2(_01876_),
    .B1(_01879_),
    .B2(_01883_),
    .C(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07141_ (.A1(net227),
    .A2(_01875_),
    .B(_01885_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07142_ (.A1(_01857_),
    .A2(_01886_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07143_ (.I(\wb_counter[12] ),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07144_ (.A1(net117),
    .A2(_01877_),
    .B(_01878_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07145_ (.I(\as2650.debug_psu[4] ),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07146_ (.I(_01747_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07147_ (.A1(_01880_),
    .A2(_01889_),
    .B(_01890_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07148_ (.A1(_01858_),
    .A2(_01887_),
    .B1(_01888_),
    .B2(_01891_),
    .C(_01884_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07149_ (.A1(net228),
    .A2(_01875_),
    .B(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07150_ (.A1(_01857_),
    .A2(_01893_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07151_ (.I(_01779_),
    .Z(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07152_ (.I(\wb_counter[13] ),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07153_ (.A1(net118),
    .A2(_01877_),
    .B(_01878_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07154_ (.I(\as2650.debug_psu[5] ),
    .Z(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07155_ (.A1(_01880_),
    .A2(_01897_),
    .B(_01890_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07156_ (.A1(_01813_),
    .A2(_01895_),
    .B1(_01896_),
    .B2(_01898_),
    .C(_01884_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07157_ (.A1(net229),
    .A2(_01875_),
    .B(_01899_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07158_ (.A1(_01894_),
    .A2(_01900_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07159_ (.I(\wb_counter[14] ),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07160_ (.A1(net119),
    .A2(_01877_),
    .B(_01878_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07161_ (.I(net173),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07162_ (.A1(_01880_),
    .A2(_01903_),
    .B(_01890_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07163_ (.A1(_01813_),
    .A2(_01901_),
    .B1(_01902_),
    .B2(_01904_),
    .C(_01884_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07164_ (.A1(net230),
    .A2(_01875_),
    .B(_01905_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07165_ (.A1(_01894_),
    .A2(_01906_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07166_ (.I(\wb_counter[15] ),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07167_ (.I(net382),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07168_ (.A1(net120),
    .A2(_01908_),
    .B(_01807_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07169_ (.I(\as2650.debug_psu[7] ),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07170_ (.A1(_01821_),
    .A2(_01910_),
    .B(_01890_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _07171_ (.A1(_01813_),
    .A2(_01907_),
    .B1(_01909_),
    .B2(_01911_),
    .C(_01802_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07172_ (.A1(net231),
    .A2(_01764_),
    .B(_01912_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07173_ (.A1(_01894_),
    .A2(_01913_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07174_ (.I(net232),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07175_ (.I(_01815_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07176_ (.I(_01915_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07177_ (.I(_01908_),
    .Z(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07178_ (.A1(net59),
    .A2(_01750_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07179_ (.A1(net62),
    .A2(net61),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07180_ (.A1(_01918_),
    .A2(_01919_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07181_ (.I(_01920_),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07182_ (.I(_01921_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07183_ (.A1(net98),
    .A2(_01917_),
    .B(_01922_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07184_ (.I(_01763_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07185_ (.A1(_01767_),
    .A2(\wb_counter[16] ),
    .B(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07186_ (.I(_01746_),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07187_ (.A1(_01914_),
    .A2(_01916_),
    .B1(_01923_),
    .B2(_01925_),
    .C(_01926_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07188_ (.I(net233),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07189_ (.A1(net105),
    .A2(_01917_),
    .B(_01922_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07190_ (.I(_01766_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07191_ (.A1(_01929_),
    .A2(\wb_counter[17] ),
    .B(_01924_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07192_ (.I(_01800_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07193_ (.A1(_01927_),
    .A2(_01916_),
    .B1(_01928_),
    .B2(_01930_),
    .C(_01931_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07194_ (.I(net234),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07195_ (.A1(net106),
    .A2(_01917_),
    .B(_01922_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07196_ (.A1(_01929_),
    .A2(\wb_counter[18] ),
    .B(_01924_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07197_ (.A1(_01932_),
    .A2(_01916_),
    .B1(_01933_),
    .B2(_01934_),
    .C(_01931_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07198_ (.I(net235),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07199_ (.I(net417),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07200_ (.A1(net107),
    .A2(_01917_),
    .B(_01936_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07201_ (.A1(_01929_),
    .A2(\wb_counter[19] ),
    .B(_01924_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07202_ (.A1(_01935_),
    .A2(_01916_),
    .B1(_01937_),
    .B2(_01938_),
    .C(_01931_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07203_ (.I(net237),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07204_ (.I(_01915_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07205_ (.I(_01908_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07206_ (.A1(net108),
    .A2(_01941_),
    .B(_01922_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07207_ (.I(_01763_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07208_ (.A1(_01929_),
    .A2(\wb_counter[20] ),
    .B(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07209_ (.A1(_01939_),
    .A2(_01940_),
    .B1(_01942_),
    .B2(_01944_),
    .C(_01931_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07210_ (.I(net238),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07211_ (.I(_01920_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07212_ (.A1(net109),
    .A2(_01941_),
    .B(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07213_ (.I(_01766_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07214_ (.A1(_01948_),
    .A2(\wb_counter[21] ),
    .B(_01943_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07215_ (.I(_01800_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07216_ (.A1(_01945_),
    .A2(_01940_),
    .B1(_01947_),
    .B2(_01949_),
    .C(_01950_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07217_ (.I(net239),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07218_ (.A1(net110),
    .A2(_01941_),
    .B(_01946_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07219_ (.A1(_01948_),
    .A2(\wb_counter[22] ),
    .B(_01943_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07220_ (.A1(_01951_),
    .A2(_01940_),
    .B1(_01952_),
    .B2(_01953_),
    .C(_01950_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07221_ (.I(net240),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07222_ (.A1(net111),
    .A2(_01941_),
    .B(_01946_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07223_ (.A1(_01948_),
    .A2(\wb_counter[23] ),
    .B(_01943_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07224_ (.A1(_01954_),
    .A2(_01940_),
    .B1(_01955_),
    .B2(_01956_),
    .C(_01950_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07225_ (.I(net241),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07226_ (.I(_01915_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07227_ (.I(_01908_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07228_ (.A1(net112),
    .A2(_01959_),
    .B(_01936_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07229_ (.I(_01763_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07230_ (.A1(_01948_),
    .A2(\wb_counter[24] ),
    .B(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07231_ (.A1(_01957_),
    .A2(_01958_),
    .B1(_01960_),
    .B2(_01962_),
    .C(_01950_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07232_ (.I(net242),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07233_ (.A1(net113),
    .A2(_01959_),
    .B(_01946_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07234_ (.I(_01766_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07235_ (.A1(_01965_),
    .A2(\wb_counter[25] ),
    .B(_01961_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07236_ (.I(_01800_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07237_ (.A1(_01963_),
    .A2(_01958_),
    .B1(_01964_),
    .B2(_01966_),
    .C(_01967_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07238_ (.I(net243),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07239_ (.A1(net99),
    .A2(_01959_),
    .B(_01921_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07240_ (.A1(_01965_),
    .A2(\wb_counter[26] ),
    .B(_01961_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07241_ (.A1(_01968_),
    .A2(_01958_),
    .B1(_01969_),
    .B2(_01970_),
    .C(_01967_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07242_ (.I(net244),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07243_ (.A1(net100),
    .A2(_01959_),
    .B(_01921_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07244_ (.A1(_01965_),
    .A2(\wb_counter[27] ),
    .B(_01961_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07245_ (.A1(_01971_),
    .A2(_01958_),
    .B1(_01972_),
    .B2(_01973_),
    .C(_01967_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07246_ (.I(net245),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07247_ (.I(_01915_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07248_ (.I(_01805_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07249_ (.A1(net101),
    .A2(_01976_),
    .B(_01936_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07250_ (.I(_01815_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07251_ (.A1(_01965_),
    .A2(\wb_counter[28] ),
    .B(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07252_ (.A1(_01974_),
    .A2(_01975_),
    .B1(_01977_),
    .B2(_01979_),
    .C(_01967_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07253_ (.I(net246),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07254_ (.A1(net102),
    .A2(_01976_),
    .B(_01936_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07255_ (.A1(_01774_),
    .A2(\wb_counter[29] ),
    .B(_01978_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07256_ (.A1(_01980_),
    .A2(_01975_),
    .B1(_01981_),
    .B2(_01982_),
    .C(_01826_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07257_ (.I(net248),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07258_ (.A1(net103),
    .A2(_01976_),
    .B(_01921_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07259_ (.A1(_01774_),
    .A2(\wb_counter[30] ),
    .B(_01978_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07260_ (.A1(_01983_),
    .A2(_01975_),
    .B1(_01984_),
    .B2(_01985_),
    .C(_01826_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07261_ (.I(net249),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _07262_ (.A1(net104),
    .A2(_01976_),
    .B1(_01918_),
    .B2(_00712_),
    .C(net417),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07263_ (.A1(_01774_),
    .A2(\wb_counter[31] ),
    .B(_01978_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _07264_ (.A1(_01986_),
    .A2(_01975_),
    .B1(net418),
    .B2(_01988_),
    .C(_01826_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07265_ (.A1(_01894_),
    .A2(net411),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07266_ (.A1(_01786_),
    .A2(_01751_),
    .A3(_01699_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07267_ (.I(_01989_),
    .Z(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07268_ (.A1(net337),
    .A2(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07269_ (.A1(_01768_),
    .A2(_01752_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07270_ (.I(_01992_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07271_ (.A1(wb_debug_cc),
    .A2(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07272_ (.A1(net338),
    .A2(_01994_),
    .B(_01780_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07273_ (.A1(net75),
    .A2(_01990_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07274_ (.A1(_01469_),
    .A2(_01993_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07275_ (.I(_01779_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07276_ (.A1(net387),
    .A2(_01996_),
    .B(_01997_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07277_ (.A1(net325),
    .A2(_01990_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07278_ (.A1(\web_behavior[0] ),
    .A2(_01993_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07279_ (.A1(net326),
    .A2(_01999_),
    .B(_01997_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07280_ (.A1(net321),
    .A2(_01990_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07281_ (.I(_01992_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07282_ (.A1(\web_behavior[1] ),
    .A2(_02001_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07283_ (.A1(net322),
    .A2(_02002_),
    .B(_01997_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07284_ (.A1(net329),
    .A2(_01989_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07285_ (.A1(wb_reset_override_en),
    .A2(_02001_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07286_ (.A1(net330),
    .A2(_02004_),
    .B(_01997_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07287_ (.A1(net91),
    .A2(_01989_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07288_ (.A1(wb_reset_override),
    .A2(_02001_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07289_ (.A1(net349),
    .A2(_02006_),
    .B(_01801_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07290_ (.A1(net378),
    .A2(_01992_),
    .B(_01760_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07291_ (.A1(net157),
    .A2(_01993_),
    .B(net379),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07292_ (.A1(net333),
    .A2(_01989_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07293_ (.A1(net174),
    .A2(_02001_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07294_ (.A1(net334),
    .A2(_02009_),
    .B(_01801_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07295_ (.I(_00712_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07296_ (.A1(net88),
    .A2(net401),
    .B(_01760_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07297_ (.A1(_02010_),
    .A2(net401),
    .B(_02011_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07298_ (.A1(net97),
    .A2(_01694_),
    .A3(_01777_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07299_ (.I(net368),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07300_ (.I(_02013_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07301_ (.A1(net64),
    .A2(_02013_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07302_ (.A1(\wb_counter[0] ),
    .A2(_02014_),
    .B(_02015_),
    .C(_01926_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07303_ (.A1(_01775_),
    .A2(\wb_counter[1] ),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07304_ (.A1(net75),
    .A2(_02013_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07305_ (.A1(_02014_),
    .A2(_02016_),
    .B(_02017_),
    .C(_01926_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07306_ (.A1(\wb_counter[0] ),
    .A2(\wb_counter[1] ),
    .A3(\wb_counter[2] ),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07307_ (.A1(_01775_),
    .A2(_01788_),
    .B(_01797_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07308_ (.A1(_02018_),
    .A2(_02019_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07309_ (.A1(net86),
    .A2(_02013_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07310_ (.A1(_02014_),
    .A2(_02020_),
    .B(_02021_),
    .C(_01926_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07311_ (.I(_02012_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07312_ (.I(_02022_),
    .Z(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07313_ (.I(_02023_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07314_ (.A1(\wb_counter[3] ),
    .A2(_02018_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07315_ (.I(_02012_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07316_ (.I(_02026_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07317_ (.A1(net321),
    .A2(_02027_),
    .B(_01760_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07318_ (.A1(_02024_),
    .A2(_02025_),
    .B(_02028_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07319_ (.A1(_01804_),
    .A2(_02018_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07320_ (.A1(_01819_),
    .A2(_02029_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07321_ (.I(_01759_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07322_ (.A1(net329),
    .A2(_02027_),
    .B(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07323_ (.A1(_02024_),
    .A2(_02030_),
    .B(_02032_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07324_ (.A1(\wb_counter[4] ),
    .A2(_02029_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07325_ (.A1(_01829_),
    .A2(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07326_ (.A1(\wb_counter[4] ),
    .A2(\wb_counter[5] ),
    .A3(_02029_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07327_ (.A1(_02034_),
    .A2(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07328_ (.A1(net91),
    .A2(_02027_),
    .B(_02031_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07329_ (.A1(_02024_),
    .A2(_02036_),
    .B(_02037_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07330_ (.A1(_01835_),
    .A2(_02035_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07331_ (.A1(_01835_),
    .A2(_02035_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07332_ (.A1(_02038_),
    .A2(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07333_ (.A1(net92),
    .A2(_02027_),
    .B(_02031_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07334_ (.A1(_02024_),
    .A2(_02040_),
    .B(_02041_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07335_ (.I(_02023_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07336_ (.A1(\wb_counter[7] ),
    .A2(_02039_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07337_ (.I(_02026_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07338_ (.A1(net93),
    .A2(_02044_),
    .B(_02031_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07339_ (.A1(_02042_),
    .A2(_02043_),
    .B(_02045_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07340_ (.A1(_01841_),
    .A2(_02039_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07341_ (.A1(_01849_),
    .A2(_02046_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07342_ (.I(_01759_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07343_ (.A1(net372),
    .A2(_02044_),
    .B(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07344_ (.A1(_02042_),
    .A2(_02047_),
    .B(_02049_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07345_ (.A1(_01841_),
    .A2(_01849_),
    .A3(_02039_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07346_ (.A1(_01859_),
    .A2(_02050_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07347_ (.A1(net364),
    .A2(_02044_),
    .B(_02048_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07348_ (.A1(_02042_),
    .A2(_02051_),
    .B(net365),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07349_ (.A1(\wb_counter[9] ),
    .A2(_02050_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07350_ (.A1(\wb_counter[10] ),
    .A2(_02053_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07351_ (.A1(net360),
    .A2(_02044_),
    .B(_02048_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07352_ (.A1(_02042_),
    .A2(_02054_),
    .B(net361),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07353_ (.I(_02023_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07354_ (.A1(_01866_),
    .A2(_02053_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07355_ (.A1(_01876_),
    .A2(_02057_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07356_ (.I(_02026_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07357_ (.A1(net370),
    .A2(_02059_),
    .B(_02048_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07358_ (.A1(_02056_),
    .A2(_02058_),
    .B(_02060_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07359_ (.A1(\wb_counter[11] ),
    .A2(\wb_counter[12] ),
    .A3(_02057_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07360_ (.A1(\wb_counter[11] ),
    .A2(_02057_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07361_ (.A1(_01887_),
    .A2(_02062_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07362_ (.A1(_02061_),
    .A2(_02063_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07363_ (.I(_01759_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07364_ (.A1(net341),
    .A2(_02059_),
    .B(_02065_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07365_ (.A1(_02056_),
    .A2(_02064_),
    .B(net342),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07366_ (.A1(\wb_counter[13] ),
    .A2(_02061_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07367_ (.A1(net345),
    .A2(_02059_),
    .B(_02065_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07368_ (.A1(_02056_),
    .A2(_02067_),
    .B(net346),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07369_ (.A1(_01895_),
    .A2(_02061_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07370_ (.A1(_01901_),
    .A2(_02069_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07371_ (.A1(net356),
    .A2(_02059_),
    .B(_02065_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07372_ (.A1(_02056_),
    .A2(_02070_),
    .B(net357),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07373_ (.I(_02012_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07374_ (.I(_02072_),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07375_ (.A1(\wb_counter[14] ),
    .A2(\wb_counter[15] ),
    .A3(_02069_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07376_ (.A1(\wb_counter[14] ),
    .A2(_02069_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07377_ (.A1(_01907_),
    .A2(_02075_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07378_ (.A1(_02074_),
    .A2(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07379_ (.I(_02026_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07380_ (.A1(net352),
    .A2(_02078_),
    .B(_02065_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07381_ (.A1(_02073_),
    .A2(_02077_),
    .B(net353),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07382_ (.A1(\wb_counter[16] ),
    .A2(_02074_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07383_ (.I(_01758_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07384_ (.I(_02081_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07385_ (.A1(net71),
    .A2(_02078_),
    .B(_02082_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07386_ (.A1(_02073_),
    .A2(_02080_),
    .B(_02083_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07387_ (.I(\wb_counter[16] ),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07388_ (.A1(_02084_),
    .A2(_02074_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07389_ (.A1(\wb_counter[17] ),
    .A2(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07390_ (.A1(net72),
    .A2(_02078_),
    .B(_02082_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07391_ (.A1(_02073_),
    .A2(_02086_),
    .B(_02087_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07392_ (.A1(\wb_counter[17] ),
    .A2(_02085_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07393_ (.A1(\wb_counter[18] ),
    .A2(_02088_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07394_ (.A1(net73),
    .A2(_02078_),
    .B(_02082_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07395_ (.A1(_02073_),
    .A2(_02089_),
    .B(_02090_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07396_ (.I(_02072_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07397_ (.A1(\wb_counter[17] ),
    .A2(\wb_counter[18] ),
    .A3(_02085_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07398_ (.A1(\wb_counter[19] ),
    .A2(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07399_ (.I(_02022_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07400_ (.A1(net74),
    .A2(_02094_),
    .B(_02082_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07401_ (.A1(_02091_),
    .A2(_02093_),
    .B(_02095_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07402_ (.I(\wb_counter[19] ),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07403_ (.A1(_02096_),
    .A2(_02092_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07404_ (.A1(\wb_counter[20] ),
    .A2(_02097_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07405_ (.I(_02081_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07406_ (.A1(net76),
    .A2(_02094_),
    .B(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07407_ (.A1(_02091_),
    .A2(_02098_),
    .B(_02100_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07408_ (.A1(\wb_counter[20] ),
    .A2(_02097_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07409_ (.A1(\wb_counter[21] ),
    .A2(_02101_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07410_ (.A1(net77),
    .A2(_02094_),
    .B(_02099_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07411_ (.A1(_02091_),
    .A2(_02102_),
    .B(_02103_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07412_ (.A1(\wb_counter[20] ),
    .A2(\wb_counter[21] ),
    .A3(_02097_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07413_ (.A1(\wb_counter[22] ),
    .A2(_02104_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07414_ (.A1(net78),
    .A2(_02094_),
    .B(_02099_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07415_ (.A1(_02091_),
    .A2(_02105_),
    .B(_02106_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07416_ (.I(_02072_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07417_ (.I(\wb_counter[22] ),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07418_ (.A1(_02108_),
    .A2(_02104_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07419_ (.A1(\wb_counter[23] ),
    .A2(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07420_ (.I(_02022_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07421_ (.A1(net79),
    .A2(_02111_),
    .B(_02099_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07422_ (.A1(_02107_),
    .A2(_02110_),
    .B(_02112_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07423_ (.A1(\wb_counter[23] ),
    .A2(_02109_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07424_ (.A1(\wb_counter[24] ),
    .A2(_02113_),
    .Z(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07425_ (.I(_02081_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07426_ (.A1(net80),
    .A2(_02111_),
    .B(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07427_ (.A1(_02107_),
    .A2(_02114_),
    .B(_02116_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07428_ (.A1(\wb_counter[23] ),
    .A2(\wb_counter[24] ),
    .A3(_02109_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07429_ (.A1(\wb_counter[25] ),
    .A2(_02117_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07430_ (.A1(net81),
    .A2(_02111_),
    .B(_02115_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07431_ (.A1(_02107_),
    .A2(_02118_),
    .B(_02119_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07432_ (.I(\wb_counter[25] ),
    .ZN(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07433_ (.A1(_02120_),
    .A2(_02117_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07434_ (.A1(\wb_counter[26] ),
    .A2(_02121_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07435_ (.A1(net82),
    .A2(_02111_),
    .B(_02115_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07436_ (.A1(_02107_),
    .A2(_02122_),
    .B(_02123_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07437_ (.I(_02072_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07438_ (.A1(\wb_counter[26] ),
    .A2(_02121_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07439_ (.A1(\wb_counter[27] ),
    .A2(_02125_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07440_ (.I(_02022_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07441_ (.A1(net83),
    .A2(_02127_),
    .B(_02115_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07442_ (.A1(_02124_),
    .A2(_02126_),
    .B(_02128_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07443_ (.A1(\wb_counter[26] ),
    .A2(\wb_counter[27] ),
    .A3(_02121_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07444_ (.A1(\wb_counter[28] ),
    .A2(_02129_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07445_ (.I(_02081_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07446_ (.A1(net84),
    .A2(_02127_),
    .B(_02131_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07447_ (.A1(_02124_),
    .A2(_02130_),
    .B(_02132_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07448_ (.I(\wb_counter[28] ),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07449_ (.A1(_02133_),
    .A2(_02129_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07450_ (.A1(\wb_counter[29] ),
    .A2(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07451_ (.A1(net85),
    .A2(_02127_),
    .B(_02131_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07452_ (.A1(_02124_),
    .A2(_02135_),
    .B(_02136_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07453_ (.A1(\wb_counter[29] ),
    .A2(_02134_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07454_ (.A1(\wb_counter[30] ),
    .A2(_02137_),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07455_ (.A1(net87),
    .A2(_02127_),
    .B(_02131_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07456_ (.A1(_02124_),
    .A2(_02138_),
    .B(_02139_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07457_ (.A1(\wb_counter[29] ),
    .A2(\wb_counter[30] ),
    .A3(_02134_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07458_ (.A1(\wb_counter[31] ),
    .A2(_02140_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07459_ (.A1(net88),
    .A2(_02023_),
    .B(_02131_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07460_ (.A1(_02014_),
    .A2(_02141_),
    .B(_02142_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07461_ (.A1(_01370_),
    .A2(_01403_),
    .A3(_01250_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07462_ (.I(_02143_),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07463_ (.A1(_00747_),
    .A2(_01683_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07464_ (.A1(_02144_),
    .A2(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07465_ (.I(_00682_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07466_ (.A1(_02147_),
    .A2(_00664_),
    .A3(_01250_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07467_ (.A1(_01425_),
    .A2(_01380_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07468_ (.A1(_01685_),
    .A2(_02149_),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07469_ (.A1(_02150_),
    .A2(_01670_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07470_ (.A1(_01673_),
    .A2(_02151_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07471_ (.I(_02147_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07472_ (.I(_01220_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07473_ (.A1(_02153_),
    .A2(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07474_ (.A1(_02148_),
    .A2(_02152_),
    .B(_02155_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07475_ (.A1(_02156_),
    .A2(_02146_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07476_ (.A1(_01407_),
    .A2(_01409_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07477_ (.I(_02158_),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07478_ (.I(_01411_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07479_ (.A1(_01409_),
    .A2(_01408_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07480_ (.I(_02161_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07481_ (.I(_02162_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07482_ (.A1(_01377_),
    .A2(_02161_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07483_ (.A1(_00928_),
    .A2(_02163_),
    .B1(_02164_),
    .B2(_00934_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07484_ (.A1(_02160_),
    .A2(_00923_),
    .A3(_02163_),
    .B(_02165_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07485_ (.A1(_01410_),
    .A2(_02161_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07486_ (.I(_02167_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07487_ (.A1(_00933_),
    .A2(_00982_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _07488_ (.A1(_00984_),
    .A2(_02163_),
    .B1(_02168_),
    .B2(_00988_),
    .C1(_02164_),
    .C2(_02169_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07489_ (.I(_02170_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07490_ (.I(_01089_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07491_ (.I(_01410_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07492_ (.A1(_01396_),
    .A2(_01419_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07493_ (.A1(_02173_),
    .A2(_02174_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07494_ (.A1(_01088_),
    .A2(_01090_),
    .A3(_02175_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07495_ (.A1(_02172_),
    .A2(_02163_),
    .B1(_02168_),
    .B2(_01629_),
    .C(_02176_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07496_ (.A1(_01601_),
    .A2(_01050_),
    .B(_01071_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07497_ (.A1(_02178_),
    .A2(_02175_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07498_ (.A1(_01601_),
    .A2(_02162_),
    .B1(_02168_),
    .B2(_01078_),
    .C(_02179_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07499_ (.A1(_01102_),
    .A2(_02175_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07500_ (.A1(_01611_),
    .A2(_02162_),
    .B1(_02168_),
    .B2(_01105_),
    .C(_02181_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07501_ (.A1(_01050_),
    .A2(_01052_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07502_ (.A1(_01056_),
    .A2(_01058_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07503_ (.A1(_01053_),
    .A2(_02162_),
    .B1(_02167_),
    .B2(_02184_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07504_ (.A1(_02183_),
    .A2(_02175_),
    .B(_02185_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07505_ (.I(_01009_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07506_ (.A1(_02187_),
    .A2(_02161_),
    .B(_02164_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07507_ (.A1(_01028_),
    .A2(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07508_ (.A1(_01057_),
    .A2(_02174_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07509_ (.A1(_02186_),
    .A2(_02189_),
    .A3(_02190_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07510_ (.A1(_02177_),
    .A2(_02180_),
    .A3(_02182_),
    .A4(_02191_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07511_ (.A1(_02166_),
    .A2(_02171_),
    .A3(_02192_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07512_ (.A1(_02159_),
    .A2(_02193_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07513_ (.I(_01001_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07514_ (.A1(\as2650.debug_psl[6] ),
    .A2(_02195_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07515_ (.I(_00789_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07516_ (.A1(\as2650.debug_psl[7] ),
    .A2(_02197_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07517_ (.A1(_02196_),
    .A2(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07518_ (.A1(_01371_),
    .A2(_02158_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07519_ (.A1(_01423_),
    .A2(_01671_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07520_ (.A1(_00750_),
    .A2(_02201_),
    .A3(_01520_),
    .A4(_02200_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07521_ (.I(_02202_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07522_ (.I(_02203_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07523_ (.I(_00708_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _07524_ (.A1(_02205_),
    .A2(_00747_),
    .A3(_01521_),
    .A4(_01668_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07525_ (.A1(_01220_),
    .A2(_02204_),
    .A3(_02206_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07526_ (.A1(_02196_),
    .A2(_02198_),
    .B(_01521_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07527_ (.A1(_01457_),
    .A2(_02159_),
    .A3(_02208_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _07528_ (.A1(_02199_),
    .A2(_02200_),
    .B(_02207_),
    .C(_02209_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07529_ (.A1(_02194_),
    .A2(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07530_ (.I(_02211_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07531_ (.I(_01396_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07532_ (.I(_01377_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07533_ (.I(_02214_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07534_ (.A1(_02213_),
    .A2(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07535_ (.A1(_02147_),
    .A2(_02154_),
    .B1(_01419_),
    .B2(_02216_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07536_ (.A1(_02212_),
    .A2(_02217_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07537_ (.A1(_01361_),
    .A2(_01364_),
    .A3(_02157_),
    .A4(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07538_ (.I(_02219_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07539_ (.I(_02220_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07540_ (.I(_02221_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07541_ (.I(\as2650.PC[0] ),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07542_ (.I(_00679_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07543_ (.A1(_02223_),
    .A2(_02224_),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07544_ (.I(\as2650.debug_psl[0] ),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07545_ (.I(_02226_),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07546_ (.I(_02227_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07547_ (.I(_01519_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07548_ (.I(_02229_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07549_ (.I(_01416_),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07550_ (.I(_01526_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07551_ (.A1(_02231_),
    .A2(_02232_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07552_ (.A1(_00739_),
    .A2(_01665_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07553_ (.A1(_01364_),
    .A2(_02234_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07554_ (.I(_02235_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07555_ (.I(_02236_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07556_ (.A1(_02230_),
    .A2(_02233_),
    .A3(_02237_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07557_ (.I(_02238_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07558_ (.I(_02239_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07559_ (.I(_02238_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07560_ (.A1(_01558_),
    .A2(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07561_ (.I(_02221_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07562_ (.A1(_02228_),
    .A2(_02240_),
    .B(_02242_),
    .C(_02243_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07563_ (.A1(_02222_),
    .A2(_02225_),
    .B(_02244_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07564_ (.I(_02245_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07565_ (.I(_01868_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07566_ (.I(_02247_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07567_ (.I(_02248_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07568_ (.I(\as2650.debug_psu[0] ),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07569_ (.I(_02250_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07570_ (.I(\as2650.debug_psu[1] ),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07571_ (.I(_02252_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07572_ (.A1(_02251_),
    .A2(_02253_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07573_ (.I(_02254_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07574_ (.I(_02255_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07575_ (.I(_02256_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07576_ (.I(_02257_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07577_ (.I(_02258_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07578_ (.I(_02259_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07579_ (.A1(_02231_),
    .A2(_02232_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07580_ (.A1(_01445_),
    .A2(_01529_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07581_ (.I(_02262_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07582_ (.I(_02263_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07583_ (.A1(_02261_),
    .A2(_02264_),
    .B(_02220_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07584_ (.I(_02265_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _07585_ (.I(_02266_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07586_ (.A1(_02249_),
    .A2(_01882_),
    .A3(_02260_),
    .A4(_02267_),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07587_ (.I(_02268_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07588_ (.I0(_02246_),
    .I1(\as2650.stack[11][0] ),
    .S(_02269_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07589_ (.I(_02270_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07590_ (.I(\as2650.debug_psl[1] ),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07591_ (.I(_02271_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07592_ (.I(_02241_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07593_ (.I(_01334_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07594_ (.I(_02239_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07595_ (.A1(_02274_),
    .A2(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07596_ (.I(_02221_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07597_ (.A1(_02272_),
    .A2(_02273_),
    .B(_02276_),
    .C(_02277_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07598_ (.I(\as2650.PC[1] ),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07599_ (.I(_02279_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07600_ (.A1(_01170_),
    .A2(_02154_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07601_ (.I(_02281_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07602_ (.I(_02282_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07603_ (.I(_02219_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07604_ (.I(_02284_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07605_ (.I(_02281_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07606_ (.A1(_00957_),
    .A2(_02279_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07607_ (.I(_02287_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07608_ (.A1(_02286_),
    .A2(_02288_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07609_ (.A1(_02280_),
    .A2(_02283_),
    .B(_02285_),
    .C(_02289_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07610_ (.A1(_02278_),
    .A2(_02290_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07611_ (.I(_02291_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07612_ (.I0(_02292_),
    .I1(\as2650.stack[11][1] ),
    .S(_02269_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07613_ (.I(_02293_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07614_ (.I(_02241_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07615_ (.A1(_01594_),
    .A2(_02275_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07616_ (.A1(\as2650.debug_psl[2] ),
    .A2(_02294_),
    .B(_02295_),
    .C(_02277_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07617_ (.I(\as2650.PC[2] ),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07618_ (.I(_02297_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07619_ (.A1(\as2650.PC[0] ),
    .A2(_02279_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07620_ (.A1(_02297_),
    .A2(_02299_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07621_ (.A1(_02286_),
    .A2(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07622_ (.A1(_02298_),
    .A2(_02283_),
    .B(_02285_),
    .C(_02301_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07623_ (.A1(_02296_),
    .A2(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07624_ (.I(_02303_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07625_ (.I0(_02304_),
    .I1(\as2650.stack[11][2] ),
    .S(_02269_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07626_ (.I(_02305_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07627_ (.I0(_01812_),
    .I1(net206),
    .S(_02239_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07628_ (.A1(\as2650.PC[0] ),
    .A2(_02279_),
    .A3(\as2650.PC[2] ),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07629_ (.A1(_00951_),
    .A2(_02307_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07630_ (.I(_02308_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07631_ (.A1(_02282_),
    .A2(_02309_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07632_ (.A1(_00951_),
    .A2(_02286_),
    .B(_02310_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07633_ (.I(_02284_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07634_ (.I0(_02306_),
    .I1(_02311_),
    .S(_02312_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07635_ (.I(_02313_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07636_ (.I0(_02314_),
    .I1(\as2650.stack[11][3] ),
    .S(_02269_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07637_ (.I(_02315_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07638_ (.I(_01615_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07639_ (.I(_02238_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07640_ (.A1(_02316_),
    .A2(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07641_ (.A1(_01492_),
    .A2(_02294_),
    .B(_02318_),
    .C(_02277_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07642_ (.I(\as2650.PC[4] ),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07643_ (.I(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07644_ (.I(_00679_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07645_ (.A1(_00951_),
    .A2(_02307_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07646_ (.A1(_02320_),
    .A2(_02323_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07647_ (.I(_02324_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07648_ (.I(_02325_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07649_ (.A1(_02322_),
    .A2(_02326_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07650_ (.A1(_02321_),
    .A2(_02283_),
    .B(_02285_),
    .C(_02327_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07651_ (.A1(_02319_),
    .A2(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07652_ (.I(_02329_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07653_ (.I(_02268_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07654_ (.I0(_02330_),
    .I1(\as2650.stack[11][4] ),
    .S(_02331_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07655_ (.I(_02332_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07656_ (.I(_01632_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07657_ (.A1(_02333_),
    .A2(_02317_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07658_ (.A1(_01486_),
    .A2(_02294_),
    .B(_02334_),
    .C(_02277_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07659_ (.I(\as2650.PC[5] ),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07660_ (.I(_02336_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07661_ (.I(_02284_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07662_ (.A1(_02320_),
    .A2(_02323_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07663_ (.A1(_02336_),
    .A2(_02339_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07664_ (.I(_02340_),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07665_ (.I(_02341_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07666_ (.A1(_02322_),
    .A2(_02342_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07667_ (.A1(_02337_),
    .A2(_02283_),
    .B(_02338_),
    .C(_02343_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07668_ (.A1(_02335_),
    .A2(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07669_ (.I(_02345_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07670_ (.I0(_02346_),
    .I1(\as2650.stack[11][5] ),
    .S(_02331_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07671_ (.I(_02347_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07672_ (.I(_00637_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07673_ (.A1(_02348_),
    .A2(_02317_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07674_ (.I(_02221_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07675_ (.A1(_01473_),
    .A2(_02294_),
    .B(_02349_),
    .C(_02350_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07676_ (.I(\as2650.PC[6] ),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07677_ (.I(_02352_),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07678_ (.I(_02282_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07679_ (.A1(_02336_),
    .A2(_02339_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07680_ (.A1(_02352_),
    .A2(_02355_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07681_ (.I(_02356_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07682_ (.A1(_02322_),
    .A2(_02357_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07683_ (.A1(_02353_),
    .A2(_02354_),
    .B(_02338_),
    .C(_02358_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07684_ (.A1(_02351_),
    .A2(_02359_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07685_ (.I(_02360_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07686_ (.I0(_02361_),
    .I1(\as2650.stack[11][6] ),
    .S(_02331_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07687_ (.I(_02362_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07688_ (.I(_02239_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07689_ (.I(_01653_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07690_ (.A1(_02364_),
    .A2(_02317_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07691_ (.A1(_01480_),
    .A2(_02363_),
    .B(_02365_),
    .C(_02350_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07692_ (.I(\as2650.PC[7] ),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07693_ (.A1(_02336_),
    .A2(_02352_),
    .A3(_02339_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07694_ (.A1(_02367_),
    .A2(_02368_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07695_ (.A1(_02282_),
    .A2(_02369_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07696_ (.A1(_02367_),
    .A2(_02354_),
    .B(_02338_),
    .C(_02370_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07697_ (.A1(_02366_),
    .A2(_02371_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07698_ (.I(_02372_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07699_ (.I0(_02373_),
    .I1(\as2650.stack[11][7] ),
    .S(_02331_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07700_ (.I(_02374_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07701_ (.I(net211),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07702_ (.I(_02238_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07703_ (.A1(_02375_),
    .A2(_02376_),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07704_ (.A1(_01851_),
    .A2(_02363_),
    .B(_02377_),
    .C(_02350_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07705_ (.I(_02224_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07706_ (.I(\as2650.PC[8] ),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07707_ (.I(\as2650.PC[7] ),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07708_ (.A1(_02381_),
    .A2(_02368_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07709_ (.A1(_02380_),
    .A2(_02382_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07710_ (.I(_02383_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07711_ (.I(_02380_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07712_ (.A1(_02385_),
    .A2(_02379_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07713_ (.I(_02312_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07714_ (.A1(_02379_),
    .A2(_02384_),
    .B(_02386_),
    .C(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07715_ (.A1(_02378_),
    .A2(_02388_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07716_ (.I(_02389_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07717_ (.I(_02268_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07718_ (.I0(_02390_),
    .I1(\as2650.stack[11][8] ),
    .S(_02391_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07719_ (.I(_02392_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07720_ (.I(_00618_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07721_ (.A1(_02393_),
    .A2(_02376_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07722_ (.A1(_01862_),
    .A2(_02363_),
    .B(_02394_),
    .C(_02350_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07723_ (.I(\as2650.PC[9] ),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07724_ (.A1(\as2650.PC[8] ),
    .A2(_02382_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _07725_ (.A1(\as2650.PC[9] ),
    .A2(_02397_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07726_ (.I(_02398_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07727_ (.A1(_02322_),
    .A2(_02399_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07728_ (.A1(_02396_),
    .A2(_02354_),
    .B(_02338_),
    .C(_02400_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07729_ (.A1(_02401_),
    .A2(_02395_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07730_ (.I(_02402_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07731_ (.I0(_02403_),
    .I1(\as2650.stack[11][9] ),
    .S(_02391_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07732_ (.I(_02404_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07733_ (.I(_01870_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07734_ (.I(net181),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07735_ (.A1(_02406_),
    .A2(_02376_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07736_ (.A1(_02405_),
    .A2(_02363_),
    .B(_02407_),
    .C(_02243_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07737_ (.I(\as2650.PC[10] ),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07738_ (.I(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07739_ (.A1(\as2650.PC[8] ),
    .A2(_02396_),
    .A3(_02382_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07740_ (.A1(_02410_),
    .A2(_02411_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07741_ (.I(_02412_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07742_ (.I(_02413_),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07743_ (.A1(_02410_),
    .A2(_02379_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07744_ (.A1(_02379_),
    .A2(_02414_),
    .B(_02415_),
    .C(_02285_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07745_ (.A1(_02416_),
    .A2(_02408_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07746_ (.I(_02417_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07747_ (.I0(_02418_),
    .I1(\as2650.stack[11][10] ),
    .S(_02391_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07748_ (.I(_02419_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07749_ (.I(_01881_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07750_ (.I(_00607_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07751_ (.A1(_02421_),
    .A2(_02376_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07752_ (.A1(_02420_),
    .A2(_02240_),
    .B(_02422_),
    .C(_02243_),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07753_ (.I(\as2650.PC[11] ),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07754_ (.A1(_02410_),
    .A2(_02411_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07755_ (.A1(_02424_),
    .A2(_02425_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07756_ (.I(_02426_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07757_ (.A1(_02224_),
    .A2(_02427_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07758_ (.A1(_02424_),
    .A2(_02354_),
    .B(_02312_),
    .C(_02428_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07759_ (.A1(_02429_),
    .A2(_02423_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07760_ (.I(_02430_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07761_ (.I0(_02431_),
    .I1(\as2650.stack[11][11] ),
    .S(_02391_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07762_ (.I(_02432_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _07763_ (.I(_00600_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07764_ (.A1(_02433_),
    .A2(_02241_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07765_ (.A1(\as2650.debug_psu[4] ),
    .A2(_02240_),
    .B(_02434_),
    .C(_02243_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07766_ (.I(\as2650.PC[12] ),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07767_ (.A1(\as2650.PC[11] ),
    .A2(_02425_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07768_ (.A1(\as2650.PC[12] ),
    .A2(_02437_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07769_ (.I(_02438_),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07770_ (.A1(_02224_),
    .A2(_02439_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07771_ (.A1(_02436_),
    .A2(_02286_),
    .B(_02312_),
    .C(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07772_ (.A1(_02435_),
    .A2(_02441_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07773_ (.I(_02442_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07774_ (.I(_02268_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07775_ (.I0(_02443_),
    .I1(\as2650.stack[11][12] ),
    .S(_02444_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07776_ (.I(_02445_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07777_ (.I(\as2650.page_reg[0] ),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07778_ (.A1(_02446_),
    .A2(_02387_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _07779_ (.I(_00594_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07780_ (.A1(_02448_),
    .A2(_02240_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07781_ (.A1(_01897_),
    .A2(_02273_),
    .B(_02449_),
    .C(_02222_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07782_ (.A1(_02447_),
    .A2(_02450_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07783_ (.I(_02451_),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07784_ (.I0(_02452_),
    .I1(\as2650.stack[11][13] ),
    .S(_02444_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07785_ (.I(_02453_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07786_ (.I(\as2650.page_reg[1] ),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07787_ (.A1(_02454_),
    .A2(_02387_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _07788_ (.I(_00590_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07789_ (.A1(_02456_),
    .A2(_02275_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07790_ (.A1(_01903_),
    .A2(_02273_),
    .B(_02457_),
    .C(_02222_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07791_ (.A1(_02455_),
    .A2(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07792_ (.I(_02459_),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07793_ (.I0(_02460_),
    .I1(\as2650.stack[11][14] ),
    .S(_02444_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07794_ (.I(_02461_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07795_ (.I(\as2650.page_reg[2] ),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07796_ (.A1(_02462_),
    .A2(_02387_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _07797_ (.I(_00584_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07798_ (.A1(_02464_),
    .A2(_02275_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07799_ (.A1(_01910_),
    .A2(_02273_),
    .B(_02465_),
    .C(_02222_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07800_ (.A1(_02463_),
    .A2(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07801_ (.I(_02467_),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07802_ (.I0(_02468_),
    .I1(\as2650.stack[11][15] ),
    .S(_02444_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07803_ (.I(_02469_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07804_ (.A1(_01851_),
    .A2(_02252_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07805_ (.I(_02470_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07806_ (.I(_02471_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07807_ (.I(_02472_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07808_ (.I(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07809_ (.I(_02474_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07810_ (.I(_02475_),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07811_ (.I(_01881_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07812_ (.I(_02233_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07813_ (.A1(_02478_),
    .A2(_02237_),
    .B(_02284_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07814_ (.A1(_01870_),
    .A2(_02477_),
    .A3(_02479_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07815_ (.A1(_02476_),
    .A2(_02480_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07816_ (.I(_02481_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07817_ (.I0(_02246_),
    .I1(\as2650.stack[2][0] ),
    .S(_02482_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07818_ (.I(_02483_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07819_ (.I0(_02292_),
    .I1(\as2650.stack[2][1] ),
    .S(_02482_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07820_ (.I(_02484_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07821_ (.I0(_02304_),
    .I1(\as2650.stack[2][2] ),
    .S(_02482_),
    .Z(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07822_ (.I(_02485_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07823_ (.I0(_02314_),
    .I1(\as2650.stack[2][3] ),
    .S(_02482_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07824_ (.I(_02486_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07825_ (.I(_02481_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07826_ (.I0(_02330_),
    .I1(\as2650.stack[2][4] ),
    .S(_02487_),
    .Z(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07827_ (.I(_02488_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07828_ (.I0(_02346_),
    .I1(\as2650.stack[2][5] ),
    .S(_02487_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07829_ (.I(_02489_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07830_ (.I0(_02361_),
    .I1(\as2650.stack[2][6] ),
    .S(_02487_),
    .Z(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07831_ (.I(_02490_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07832_ (.I0(_02373_),
    .I1(\as2650.stack[2][7] ),
    .S(_02487_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07833_ (.I(_02491_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07834_ (.I(_02481_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07835_ (.I0(_02390_),
    .I1(\as2650.stack[2][8] ),
    .S(_02492_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07836_ (.I(_02493_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07837_ (.I0(_02403_),
    .I1(\as2650.stack[2][9] ),
    .S(_02492_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07838_ (.I(_02494_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07839_ (.I0(_02418_),
    .I1(\as2650.stack[2][10] ),
    .S(_02492_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07840_ (.I(_02495_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07841_ (.I0(_02431_),
    .I1(\as2650.stack[2][11] ),
    .S(_02492_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07842_ (.I(_02496_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07843_ (.I(_02481_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07844_ (.I0(_02443_),
    .I1(\as2650.stack[2][12] ),
    .S(_02497_),
    .Z(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07845_ (.I(_02498_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07846_ (.I0(_02452_),
    .I1(\as2650.stack[2][13] ),
    .S(_02497_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07847_ (.I(_02499_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07848_ (.I0(_02460_),
    .I1(\as2650.stack[2][14] ),
    .S(_02497_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07849_ (.I(_02500_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07850_ (.I0(_02468_),
    .I1(\as2650.stack[2][15] ),
    .S(_02497_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07851_ (.I(_02501_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07852_ (.A1(_02260_),
    .A2(_02480_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07853_ (.I(_02502_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07854_ (.I0(_02246_),
    .I1(\as2650.stack[3][0] ),
    .S(_02503_),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07855_ (.I(_02504_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07856_ (.I0(_02292_),
    .I1(\as2650.stack[3][1] ),
    .S(_02503_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07857_ (.I(_02505_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07858_ (.I0(_02304_),
    .I1(\as2650.stack[3][2] ),
    .S(_02503_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07859_ (.I(_02506_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07860_ (.I0(_02314_),
    .I1(\as2650.stack[3][3] ),
    .S(_02503_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07861_ (.I(_02507_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07862_ (.I(_02502_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07863_ (.I0(_02330_),
    .I1(\as2650.stack[3][4] ),
    .S(_02508_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07864_ (.I(_02509_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07865_ (.I0(_02346_),
    .I1(\as2650.stack[3][5] ),
    .S(_02508_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07866_ (.I(_02510_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07867_ (.I0(_02361_),
    .I1(\as2650.stack[3][6] ),
    .S(_02508_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07868_ (.I(_02511_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07869_ (.I0(_02373_),
    .I1(\as2650.stack[3][7] ),
    .S(_02508_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07870_ (.I(_02512_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07871_ (.I(_02502_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07872_ (.I0(_02390_),
    .I1(\as2650.stack[3][8] ),
    .S(_02513_),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07873_ (.I(_02514_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07874_ (.I0(_02403_),
    .I1(\as2650.stack[3][9] ),
    .S(_02513_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07875_ (.I(_02515_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07876_ (.I0(_02418_),
    .I1(\as2650.stack[3][10] ),
    .S(_02513_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07877_ (.I(_02516_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07878_ (.I0(_02431_),
    .I1(\as2650.stack[3][11] ),
    .S(_02513_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07879_ (.I(_02517_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07880_ (.I(_02502_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07881_ (.I0(_02443_),
    .I1(\as2650.stack[3][12] ),
    .S(_02518_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07882_ (.I(_02519_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07883_ (.I0(_02452_),
    .I1(\as2650.stack[3][13] ),
    .S(_02518_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07884_ (.I(_02520_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07885_ (.I0(_02460_),
    .I1(\as2650.stack[3][14] ),
    .S(_02518_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07886_ (.I(_02521_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07887_ (.I0(_02468_),
    .I1(\as2650.stack[3][15] ),
    .S(_02518_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07888_ (.I(_02522_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07889_ (.I(\as2650.debug_psu[3] ),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07890_ (.I(_02523_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07891_ (.A1(_02250_),
    .A2(_02252_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07892_ (.A1(\as2650.debug_psu[2] ),
    .A2(_02525_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07893_ (.A1(_02524_),
    .A2(_02267_),
    .A3(_02526_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07894_ (.I(_02527_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07895_ (.I0(_02246_),
    .I1(\as2650.stack[0][0] ),
    .S(_02528_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07896_ (.I(_02529_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07897_ (.I0(_02292_),
    .I1(\as2650.stack[0][1] ),
    .S(_02528_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07898_ (.I(_02530_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07899_ (.I0(_02304_),
    .I1(\as2650.stack[0][2] ),
    .S(_02528_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07900_ (.I(_02531_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07901_ (.I0(_02314_),
    .I1(\as2650.stack[0][3] ),
    .S(_02528_),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07902_ (.I(_02532_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07903_ (.I(_02527_),
    .Z(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07904_ (.I0(_02330_),
    .I1(\as2650.stack[0][4] ),
    .S(_02533_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07905_ (.I(_02534_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07906_ (.I0(_02346_),
    .I1(\as2650.stack[0][5] ),
    .S(_02533_),
    .Z(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07907_ (.I(_02535_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07908_ (.I0(_02361_),
    .I1(\as2650.stack[0][6] ),
    .S(_02533_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07909_ (.I(_02536_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07910_ (.I0(_02373_),
    .I1(\as2650.stack[0][7] ),
    .S(_02533_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07911_ (.I(_02537_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07912_ (.I(_02527_),
    .Z(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07913_ (.I0(_02390_),
    .I1(\as2650.stack[0][8] ),
    .S(_02538_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07914_ (.I(_02539_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07915_ (.I0(_02403_),
    .I1(\as2650.stack[0][9] ),
    .S(_02538_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07916_ (.I(_02540_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07917_ (.I0(_02418_),
    .I1(\as2650.stack[0][10] ),
    .S(_02538_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07918_ (.I(_02541_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07919_ (.I0(_02431_),
    .I1(\as2650.stack[0][11] ),
    .S(_02538_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07920_ (.I(_02542_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07921_ (.I(_02527_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07922_ (.I0(_02443_),
    .I1(\as2650.stack[0][12] ),
    .S(_02543_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07923_ (.I(_02544_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07924_ (.I0(_02452_),
    .I1(\as2650.stack[0][13] ),
    .S(_02543_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07925_ (.I(_02545_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07926_ (.I0(_02460_),
    .I1(\as2650.stack[0][14] ),
    .S(_02543_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07927_ (.I(_02546_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07928_ (.I0(_02468_),
    .I1(\as2650.stack[0][15] ),
    .S(_02543_),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07929_ (.I(_02547_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07930_ (.I(_02245_),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07931_ (.I(_02265_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _07932_ (.A1(_02405_),
    .A2(_02477_),
    .A3(_02549_),
    .A4(_02476_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07933_ (.I(_02550_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07934_ (.I0(\as2650.stack[14][0] ),
    .I1(_02548_),
    .S(_02551_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07935_ (.I(_02552_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07936_ (.I(_02291_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07937_ (.I0(\as2650.stack[14][1] ),
    .I1(_02553_),
    .S(_02551_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07938_ (.I(_02554_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07939_ (.I(_02303_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07940_ (.I0(\as2650.stack[14][2] ),
    .I1(_02555_),
    .S(_02551_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07941_ (.I(_02556_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07942_ (.I(_02313_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07943_ (.I0(\as2650.stack[14][3] ),
    .I1(_02557_),
    .S(_02551_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07944_ (.I(_02558_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07945_ (.I(_02329_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07946_ (.I(_02550_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07947_ (.I0(\as2650.stack[14][4] ),
    .I1(_02559_),
    .S(_02560_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07948_ (.I(_02561_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07949_ (.I(_02345_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07950_ (.I0(\as2650.stack[14][5] ),
    .I1(_02562_),
    .S(_02560_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07951_ (.I(_02563_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07952_ (.I(_02360_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07953_ (.I0(\as2650.stack[14][6] ),
    .I1(_02564_),
    .S(_02560_),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07954_ (.I(_02565_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07955_ (.I(_02372_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07956_ (.I0(\as2650.stack[14][7] ),
    .I1(_02566_),
    .S(_02560_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07957_ (.I(_02567_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07958_ (.I(_02389_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07959_ (.I(_02550_),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07960_ (.I0(\as2650.stack[14][8] ),
    .I1(_02568_),
    .S(_02569_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07961_ (.I(_02570_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07962_ (.I(_02402_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07963_ (.I0(\as2650.stack[14][9] ),
    .I1(_02571_),
    .S(_02569_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07964_ (.I(_02572_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07965_ (.I(_02417_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07966_ (.I0(\as2650.stack[14][10] ),
    .I1(_02573_),
    .S(_02569_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07967_ (.I(_02574_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07968_ (.I(_02430_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07969_ (.I0(\as2650.stack[14][11] ),
    .I1(_02575_),
    .S(_02569_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07970_ (.I(_02576_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07971_ (.I(_02442_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07972_ (.I(_02550_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07973_ (.I0(\as2650.stack[14][12] ),
    .I1(_02577_),
    .S(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07974_ (.I(_02579_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07975_ (.I(_02451_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07976_ (.I0(\as2650.stack[14][13] ),
    .I1(_02580_),
    .S(_02578_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07977_ (.I(_02581_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07978_ (.I(_02459_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07979_ (.I0(\as2650.stack[14][14] ),
    .I1(_02582_),
    .S(_02578_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07980_ (.I(_02583_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07981_ (.I(_02467_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07982_ (.I0(\as2650.stack[14][15] ),
    .I1(_02584_),
    .S(_02578_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07983_ (.I(_02585_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07984_ (.A1(_02251_),
    .A2(_01861_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07985_ (.I(_02586_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07986_ (.I(_02587_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07987_ (.I(_02588_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07988_ (.I(_02589_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07989_ (.I(_02590_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07990_ (.I(_02591_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _07991_ (.A1(_02405_),
    .A2(_02477_),
    .A3(_02266_),
    .A4(_02592_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07992_ (.I(_02593_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07993_ (.I0(\as2650.stack[13][0] ),
    .I1(_02548_),
    .S(_02594_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07994_ (.I(_02595_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07995_ (.I0(\as2650.stack[13][1] ),
    .I1(_02553_),
    .S(_02594_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07996_ (.I(_02596_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07997_ (.I0(\as2650.stack[13][2] ),
    .I1(_02555_),
    .S(_02594_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07998_ (.I(_02597_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07999_ (.I0(\as2650.stack[13][3] ),
    .I1(_02557_),
    .S(_02594_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08000_ (.I(_02598_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08001_ (.I(_02593_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08002_ (.I0(\as2650.stack[13][4] ),
    .I1(_02559_),
    .S(_02599_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08003_ (.I(_02600_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08004_ (.I0(\as2650.stack[13][5] ),
    .I1(_02562_),
    .S(_02599_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08005_ (.I(_02601_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08006_ (.I0(\as2650.stack[13][6] ),
    .I1(_02564_),
    .S(_02599_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08007_ (.I(_02602_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08008_ (.I0(\as2650.stack[13][7] ),
    .I1(_02566_),
    .S(_02599_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08009_ (.I(_02603_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08010_ (.I(_02593_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08011_ (.I0(\as2650.stack[13][8] ),
    .I1(_02568_),
    .S(_02604_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08012_ (.I(_02605_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08013_ (.I0(\as2650.stack[13][9] ),
    .I1(_02571_),
    .S(_02604_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08014_ (.I(_02606_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08015_ (.I0(\as2650.stack[13][10] ),
    .I1(_02573_),
    .S(_02604_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08016_ (.I(_02607_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08017_ (.I0(\as2650.stack[13][11] ),
    .I1(_02575_),
    .S(_02604_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08018_ (.I(_02608_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08019_ (.I(_02593_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08020_ (.I0(\as2650.stack[13][12] ),
    .I1(_02577_),
    .S(_02609_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08021_ (.I(_02610_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08022_ (.I0(\as2650.stack[13][13] ),
    .I1(_02580_),
    .S(_02609_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08023_ (.I(_02611_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08024_ (.I0(\as2650.stack[13][14] ),
    .I1(_02582_),
    .S(_02609_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08025_ (.I(_02612_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08026_ (.I0(\as2650.stack[13][15] ),
    .I1(_02584_),
    .S(_02609_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08027_ (.I(_02613_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08028_ (.I(_02245_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08029_ (.I(_02523_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08030_ (.A1(_02248_),
    .A2(_02615_),
    .A3(_02479_),
    .A4(_02525_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08031_ (.I(_02616_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08032_ (.I0(\as2650.stack[12][0] ),
    .I1(_02614_),
    .S(_02617_),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08033_ (.I(_02618_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08034_ (.I(_02291_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08035_ (.I0(\as2650.stack[12][1] ),
    .I1(_02619_),
    .S(_02617_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08036_ (.I(_02620_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08037_ (.I(_02303_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08038_ (.I0(\as2650.stack[12][2] ),
    .I1(_02621_),
    .S(_02617_),
    .Z(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08039_ (.I(_02622_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08040_ (.I(_02313_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08041_ (.I0(\as2650.stack[12][3] ),
    .I1(_02623_),
    .S(_02617_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08042_ (.I(_02624_),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08043_ (.I(_02329_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08044_ (.I(_02616_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08045_ (.I0(\as2650.stack[12][4] ),
    .I1(_02625_),
    .S(_02626_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08046_ (.I(_02627_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08047_ (.I(_02345_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08048_ (.I0(\as2650.stack[12][5] ),
    .I1(_02628_),
    .S(_02626_),
    .Z(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08049_ (.I(_02629_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08050_ (.I(_02360_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08051_ (.I0(\as2650.stack[12][6] ),
    .I1(_02630_),
    .S(_02626_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08052_ (.I(_02631_),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08053_ (.I(_02372_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08054_ (.I0(\as2650.stack[12][7] ),
    .I1(_02632_),
    .S(_02626_),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08055_ (.I(_02633_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08056_ (.I(_02389_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08057_ (.I(_02616_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08058_ (.I0(\as2650.stack[12][8] ),
    .I1(_02634_),
    .S(_02635_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08059_ (.I(_02636_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08060_ (.I(_02402_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08061_ (.I0(\as2650.stack[12][9] ),
    .I1(_02637_),
    .S(_02635_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08062_ (.I(_02638_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08063_ (.I(_02417_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08064_ (.I0(\as2650.stack[12][10] ),
    .I1(_02639_),
    .S(_02635_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08065_ (.I(_02640_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08066_ (.I(_02430_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08067_ (.I0(\as2650.stack[12][11] ),
    .I1(_02641_),
    .S(_02635_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08068_ (.I(_02642_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08069_ (.I(_02442_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08070_ (.I(_02616_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08071_ (.I0(\as2650.stack[12][12] ),
    .I1(_02643_),
    .S(_02644_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08072_ (.I(_02645_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08073_ (.I(_02451_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08074_ (.I0(\as2650.stack[12][13] ),
    .I1(_02646_),
    .S(_02644_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08075_ (.I(_02647_),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08076_ (.I(_02459_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08077_ (.I0(\as2650.stack[12][14] ),
    .I1(_02648_),
    .S(_02644_),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08078_ (.I(_02649_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08079_ (.I(_02467_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08080_ (.I0(\as2650.stack[12][15] ),
    .I1(_02650_),
    .S(_02644_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08081_ (.I(_02651_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08082_ (.I(_02245_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08083_ (.A1(_01882_),
    .A2(_02267_),
    .A3(_02526_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08084_ (.I(_02653_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08085_ (.I0(_02652_),
    .I1(\as2650.stack[8][0] ),
    .S(_02654_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08086_ (.I(_02655_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08087_ (.I(_02291_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08088_ (.I0(_02656_),
    .I1(\as2650.stack[8][1] ),
    .S(_02654_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08089_ (.I(_02657_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08090_ (.I(_02303_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08091_ (.I0(_02658_),
    .I1(\as2650.stack[8][2] ),
    .S(_02654_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08092_ (.I(_02659_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08093_ (.I(_02313_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08094_ (.I0(_02660_),
    .I1(\as2650.stack[8][3] ),
    .S(_02654_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08095_ (.I(_02661_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08096_ (.I(_02329_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08097_ (.I(_02653_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08098_ (.I0(_02662_),
    .I1(\as2650.stack[8][4] ),
    .S(_02663_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08099_ (.I(_02664_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08100_ (.I(_02345_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08101_ (.I0(_02665_),
    .I1(\as2650.stack[8][5] ),
    .S(_02663_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08102_ (.I(_02666_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08103_ (.I(_02360_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08104_ (.I0(_02667_),
    .I1(\as2650.stack[8][6] ),
    .S(_02663_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08105_ (.I(_02668_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08106_ (.I(_02372_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08107_ (.I0(_02669_),
    .I1(\as2650.stack[8][7] ),
    .S(_02663_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08108_ (.I(_02670_),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08109_ (.I(_02389_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08110_ (.I(_02653_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08111_ (.I0(_02671_),
    .I1(\as2650.stack[8][8] ),
    .S(_02672_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08112_ (.I(_02673_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08113_ (.I(_02402_),
    .Z(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08114_ (.I0(_02674_),
    .I1(\as2650.stack[8][9] ),
    .S(_02672_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08115_ (.I(_02675_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08116_ (.I(_02417_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08117_ (.I0(_02676_),
    .I1(\as2650.stack[8][10] ),
    .S(_02672_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08118_ (.I(_02677_),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08119_ (.I(_02430_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08120_ (.I0(_02678_),
    .I1(\as2650.stack[8][11] ),
    .S(_02672_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08121_ (.I(_02679_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08122_ (.I(_02442_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08123_ (.I(_02653_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08124_ (.I0(_02680_),
    .I1(\as2650.stack[8][12] ),
    .S(_02681_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08125_ (.I(_02682_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08126_ (.I(_02451_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08127_ (.I0(_02683_),
    .I1(\as2650.stack[8][13] ),
    .S(_02681_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08128_ (.I(_02684_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08129_ (.I(_02459_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08130_ (.I0(_02685_),
    .I1(\as2650.stack[8][14] ),
    .S(_02681_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08131_ (.I(_02686_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08132_ (.I(_02467_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08133_ (.I0(_02687_),
    .I1(\as2650.stack[8][15] ),
    .S(_02681_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08134_ (.I(_02688_),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08135_ (.A1(_01871_),
    .A2(_02524_),
    .A3(_02260_),
    .A4(_02267_),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08136_ (.I(_02689_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08137_ (.I0(_02652_),
    .I1(\as2650.stack[7][0] ),
    .S(_02690_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08138_ (.I(_02691_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08139_ (.I0(_02656_),
    .I1(\as2650.stack[7][1] ),
    .S(_02690_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08140_ (.I(_02692_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08141_ (.I0(_02658_),
    .I1(\as2650.stack[7][2] ),
    .S(_02690_),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08142_ (.I(_02693_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08143_ (.I0(_02660_),
    .I1(\as2650.stack[7][3] ),
    .S(_02690_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08144_ (.I(_02694_),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08145_ (.I(_02689_),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08146_ (.I0(_02662_),
    .I1(\as2650.stack[7][4] ),
    .S(_02695_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08147_ (.I(_02696_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08148_ (.I0(_02665_),
    .I1(\as2650.stack[7][5] ),
    .S(_02695_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08149_ (.I(_02697_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08150_ (.I0(_02667_),
    .I1(\as2650.stack[7][6] ),
    .S(_02695_),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08151_ (.I(_02698_),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08152_ (.I0(_02669_),
    .I1(\as2650.stack[7][7] ),
    .S(_02695_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08153_ (.I(_02699_),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08154_ (.I(_02689_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08155_ (.I0(_02671_),
    .I1(\as2650.stack[7][8] ),
    .S(_02700_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08156_ (.I(_02701_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08157_ (.I0(_02674_),
    .I1(\as2650.stack[7][9] ),
    .S(_02700_),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08158_ (.I(_02702_),
    .Z(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08159_ (.I0(_02676_),
    .I1(\as2650.stack[7][10] ),
    .S(_02700_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08160_ (.I(_02703_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08161_ (.I0(_02678_),
    .I1(\as2650.stack[7][11] ),
    .S(_02700_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08162_ (.I(_02704_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08163_ (.I(_02689_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08164_ (.I0(_02680_),
    .I1(\as2650.stack[7][12] ),
    .S(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08165_ (.I(_02706_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08166_ (.I0(_02683_),
    .I1(\as2650.stack[7][13] ),
    .S(_02705_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08167_ (.I(_02707_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08168_ (.I0(_02685_),
    .I1(\as2650.stack[7][14] ),
    .S(_02705_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08169_ (.I(_02708_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08170_ (.I0(_02687_),
    .I1(\as2650.stack[7][15] ),
    .S(_02705_),
    .Z(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08171_ (.I(_02709_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _08172_ (.A1(_02405_),
    .A2(_02615_),
    .A3(_02266_),
    .A4(_02476_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08173_ (.I(_02710_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08174_ (.I0(\as2650.stack[6][0] ),
    .I1(_02614_),
    .S(_02711_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08175_ (.I(_02712_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08176_ (.I0(\as2650.stack[6][1] ),
    .I1(_02619_),
    .S(_02711_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08177_ (.I(_02713_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08178_ (.I0(\as2650.stack[6][2] ),
    .I1(_02621_),
    .S(_02711_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08179_ (.I(_02714_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08180_ (.I0(\as2650.stack[6][3] ),
    .I1(_02623_),
    .S(_02711_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08181_ (.I(_02715_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08182_ (.I(_02710_),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08183_ (.I0(\as2650.stack[6][4] ),
    .I1(_02625_),
    .S(_02716_),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08184_ (.I(_02717_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08185_ (.I0(\as2650.stack[6][5] ),
    .I1(_02628_),
    .S(_02716_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08186_ (.I(_02718_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08187_ (.I0(\as2650.stack[6][6] ),
    .I1(_02630_),
    .S(_02716_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08188_ (.I(_02719_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08189_ (.I0(\as2650.stack[6][7] ),
    .I1(_02632_),
    .S(_02716_),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08190_ (.I(_02720_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08191_ (.I(_02710_),
    .Z(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08192_ (.I0(\as2650.stack[6][8] ),
    .I1(_02634_),
    .S(_02721_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08193_ (.I(_02722_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08194_ (.I0(\as2650.stack[6][9] ),
    .I1(_02637_),
    .S(_02721_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08195_ (.I(_02723_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08196_ (.I0(\as2650.stack[6][10] ),
    .I1(_02639_),
    .S(_02721_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08197_ (.I(_02724_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08198_ (.I0(\as2650.stack[6][11] ),
    .I1(_02641_),
    .S(_02721_),
    .Z(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08199_ (.I(_02725_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08200_ (.I(_02710_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08201_ (.I0(\as2650.stack[6][12] ),
    .I1(_02643_),
    .S(_02726_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08202_ (.I(_02727_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08203_ (.I0(\as2650.stack[6][13] ),
    .I1(_02646_),
    .S(_02726_),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08204_ (.I(_02728_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08205_ (.I0(\as2650.stack[6][14] ),
    .I1(_02648_),
    .S(_02726_),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08206_ (.I(_02729_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08207_ (.I0(\as2650.stack[6][15] ),
    .I1(_02650_),
    .S(_02726_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08208_ (.I(_02730_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _08209_ (.A1(_01870_),
    .A2(_02615_),
    .A3(_02266_),
    .A4(_02592_),
    .Z(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08210_ (.I(_02731_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08211_ (.I0(\as2650.stack[5][0] ),
    .I1(_02614_),
    .S(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08212_ (.I(_02733_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08213_ (.I0(\as2650.stack[5][1] ),
    .I1(_02619_),
    .S(_02732_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08214_ (.I(_02734_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08215_ (.I0(\as2650.stack[5][2] ),
    .I1(_02621_),
    .S(_02732_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08216_ (.I(_02735_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08217_ (.I0(\as2650.stack[5][3] ),
    .I1(_02623_),
    .S(_02732_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08218_ (.I(_02736_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08219_ (.I(_02731_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08220_ (.I0(\as2650.stack[5][4] ),
    .I1(_02625_),
    .S(_02737_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08221_ (.I(_02738_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08222_ (.I0(\as2650.stack[5][5] ),
    .I1(_02628_),
    .S(_02737_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08223_ (.I(_02739_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08224_ (.I0(\as2650.stack[5][6] ),
    .I1(_02630_),
    .S(_02737_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08225_ (.I(_02740_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08226_ (.I0(\as2650.stack[5][7] ),
    .I1(_02632_),
    .S(_02737_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08227_ (.I(_02741_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08228_ (.I(_02731_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08229_ (.I0(\as2650.stack[5][8] ),
    .I1(_02634_),
    .S(_02742_),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08230_ (.I(_02743_),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08231_ (.I0(\as2650.stack[5][9] ),
    .I1(_02637_),
    .S(_02742_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08232_ (.I(_02744_),
    .Z(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08233_ (.I0(\as2650.stack[5][10] ),
    .I1(_02639_),
    .S(_02742_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08234_ (.I(_02745_),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08235_ (.I0(\as2650.stack[5][11] ),
    .I1(_02641_),
    .S(_02742_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08236_ (.I(_02746_),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08237_ (.I(_02731_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08238_ (.I0(\as2650.stack[5][12] ),
    .I1(_02643_),
    .S(_02747_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08239_ (.I(_02748_),
    .Z(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08240_ (.I0(\as2650.stack[5][13] ),
    .I1(_02646_),
    .S(_02747_),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08241_ (.I(_02749_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08242_ (.I0(\as2650.stack[5][14] ),
    .I1(_02648_),
    .S(_02747_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08243_ (.I(_02750_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08244_ (.I0(\as2650.stack[5][15] ),
    .I1(_02650_),
    .S(_02747_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08245_ (.I(_02751_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08246_ (.A1(_02249_),
    .A2(_02420_),
    .A3(_02549_),
    .A4(_02476_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08247_ (.I(_02752_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08248_ (.I0(_02652_),
    .I1(\as2650.stack[10][0] ),
    .S(_02753_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08249_ (.I(_02754_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08250_ (.I0(_02656_),
    .I1(\as2650.stack[10][1] ),
    .S(_02753_),
    .Z(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08251_ (.I(_02755_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08252_ (.I0(_02658_),
    .I1(\as2650.stack[10][2] ),
    .S(_02753_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08253_ (.I(_02756_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08254_ (.I0(_02660_),
    .I1(\as2650.stack[10][3] ),
    .S(_02753_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08255_ (.I(_02757_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08256_ (.I(_02752_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08257_ (.I0(_02662_),
    .I1(\as2650.stack[10][4] ),
    .S(_02758_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08258_ (.I(_02759_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08259_ (.I0(_02665_),
    .I1(\as2650.stack[10][5] ),
    .S(_02758_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08260_ (.I(_02760_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08261_ (.I0(_02667_),
    .I1(\as2650.stack[10][6] ),
    .S(_02758_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08262_ (.I(_02761_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08263_ (.I0(_02669_),
    .I1(\as2650.stack[10][7] ),
    .S(_02758_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08264_ (.I(_02762_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08265_ (.I(_02752_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08266_ (.I0(_02671_),
    .I1(\as2650.stack[10][8] ),
    .S(_02763_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08267_ (.I(_02764_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08268_ (.I0(_02674_),
    .I1(\as2650.stack[10][9] ),
    .S(_02763_),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08269_ (.I(_02765_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08270_ (.I0(_02676_),
    .I1(\as2650.stack[10][10] ),
    .S(_02763_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08271_ (.I(_02766_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08272_ (.I0(_02678_),
    .I1(\as2650.stack[10][11] ),
    .S(_02763_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08273_ (.I(_02767_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08274_ (.I(_02752_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08275_ (.I0(_02680_),
    .I1(\as2650.stack[10][12] ),
    .S(_02768_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08276_ (.I(_02769_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08277_ (.I0(_02683_),
    .I1(\as2650.stack[10][13] ),
    .S(_02768_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08278_ (.I(_02770_),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08279_ (.I0(_02685_),
    .I1(\as2650.stack[10][14] ),
    .S(_02768_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08280_ (.I(_02771_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08281_ (.I0(_02687_),
    .I1(\as2650.stack[10][15] ),
    .S(_02768_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08282_ (.I(_02772_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08283_ (.A1(_02248_),
    .A2(_02477_),
    .A3(_02479_),
    .A4(_02525_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08284_ (.I(_02773_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08285_ (.I0(\as2650.stack[4][0] ),
    .I1(_02614_),
    .S(_02774_),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08286_ (.I(_02775_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08287_ (.I0(\as2650.stack[4][1] ),
    .I1(_02619_),
    .S(_02774_),
    .Z(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08288_ (.I(_02776_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08289_ (.I0(\as2650.stack[4][2] ),
    .I1(_02621_),
    .S(_02774_),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08290_ (.I(_02777_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08291_ (.I0(\as2650.stack[4][3] ),
    .I1(_02623_),
    .S(_02774_),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08292_ (.I(_02778_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08293_ (.I(_02773_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08294_ (.I0(\as2650.stack[4][4] ),
    .I1(_02625_),
    .S(_02779_),
    .Z(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08295_ (.I(_02780_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08296_ (.I0(\as2650.stack[4][5] ),
    .I1(_02628_),
    .S(_02779_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08297_ (.I(_02781_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08298_ (.I0(\as2650.stack[4][6] ),
    .I1(_02630_),
    .S(_02779_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08299_ (.I(_02782_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08300_ (.I0(\as2650.stack[4][7] ),
    .I1(_02632_),
    .S(_02779_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08301_ (.I(_02783_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08302_ (.I(_02773_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08303_ (.I0(\as2650.stack[4][8] ),
    .I1(_02634_),
    .S(_02784_),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08304_ (.I(_02785_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08305_ (.I0(\as2650.stack[4][9] ),
    .I1(_02637_),
    .S(_02784_),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08306_ (.I(_02786_),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08307_ (.I0(\as2650.stack[4][10] ),
    .I1(_02639_),
    .S(_02784_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08308_ (.I(_02787_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08309_ (.I0(\as2650.stack[4][11] ),
    .I1(_02641_),
    .S(_02784_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08310_ (.I(_02788_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08311_ (.I(_02773_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08312_ (.I0(\as2650.stack[4][12] ),
    .I1(_02643_),
    .S(_02789_),
    .Z(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08313_ (.I(_02790_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08314_ (.I0(\as2650.stack[4][13] ),
    .I1(_02646_),
    .S(_02789_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08315_ (.I(_02791_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08316_ (.I0(\as2650.stack[4][14] ),
    .I1(_02648_),
    .S(_02789_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08317_ (.I(_02792_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08318_ (.I0(\as2650.stack[4][15] ),
    .I1(_02650_),
    .S(_02789_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08319_ (.I(_02793_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08320_ (.A1(_01871_),
    .A2(_02420_),
    .A3(_02260_),
    .A4(_02549_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08321_ (.I(_02794_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08322_ (.I0(_02652_),
    .I1(\as2650.stack[15][0] ),
    .S(_02795_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08323_ (.I(_02796_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08324_ (.I0(_02656_),
    .I1(\as2650.stack[15][1] ),
    .S(_02795_),
    .Z(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08325_ (.I(_02797_),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08326_ (.I0(_02658_),
    .I1(\as2650.stack[15][2] ),
    .S(_02795_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08327_ (.I(_02798_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08328_ (.I0(_02660_),
    .I1(\as2650.stack[15][3] ),
    .S(_02795_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08329_ (.I(_02799_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08330_ (.I(_02794_),
    .Z(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08331_ (.I0(_02662_),
    .I1(\as2650.stack[15][4] ),
    .S(_02800_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08332_ (.I(_02801_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08333_ (.I0(_02665_),
    .I1(\as2650.stack[15][5] ),
    .S(_02800_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08334_ (.I(_02802_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08335_ (.I0(_02667_),
    .I1(\as2650.stack[15][6] ),
    .S(_02800_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08336_ (.I(_02803_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08337_ (.I0(_02669_),
    .I1(\as2650.stack[15][7] ),
    .S(_02800_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08338_ (.I(_02804_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08339_ (.I(_02794_),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08340_ (.I0(_02671_),
    .I1(\as2650.stack[15][8] ),
    .S(_02805_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08341_ (.I(_02806_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08342_ (.I0(_02674_),
    .I1(\as2650.stack[15][9] ),
    .S(_02805_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08343_ (.I(_02807_),
    .Z(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08344_ (.I0(_02676_),
    .I1(\as2650.stack[15][10] ),
    .S(_02805_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08345_ (.I(_02808_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08346_ (.I0(_02678_),
    .I1(\as2650.stack[15][11] ),
    .S(_02805_),
    .Z(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08347_ (.I(_02809_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08348_ (.I(_02794_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08349_ (.I0(_02680_),
    .I1(\as2650.stack[15][12] ),
    .S(_02810_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08350_ (.I(_02811_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08351_ (.I0(_02683_),
    .I1(\as2650.stack[15][13] ),
    .S(_02810_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08352_ (.I(_02812_),
    .Z(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08353_ (.I0(_02685_),
    .I1(\as2650.stack[15][14] ),
    .S(_02810_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08354_ (.I(_02813_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08355_ (.I0(_02687_),
    .I1(\as2650.stack[15][15] ),
    .S(_02810_),
    .Z(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08356_ (.I(_02814_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08357_ (.I(_00811_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08358_ (.I(_02815_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08359_ (.I(_02816_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08360_ (.I(_02817_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08361_ (.I(_00771_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08362_ (.I(_02819_),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08363_ (.I(_02820_),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08364_ (.I(_02821_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08365_ (.I(_02145_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08366_ (.A1(_01185_),
    .A2(_01446_),
    .A3(_02159_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08367_ (.A1(_02144_),
    .A2(_01360_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08368_ (.A1(_01675_),
    .A2(_01684_),
    .B(_02825_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _08369_ (.A1(_02823_),
    .A2(_02824_),
    .A3(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08370_ (.A1(_01423_),
    .A2(_01671_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08371_ (.I(_02828_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08372_ (.I(_02829_),
    .Z(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08373_ (.I(_02830_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08374_ (.I(_02831_),
    .Z(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08375_ (.I(_02832_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08376_ (.I(_02833_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08377_ (.A1(_02834_),
    .A2(_01427_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08378_ (.A1(_01412_),
    .A2(_01420_),
    .A3(_01672_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08379_ (.A1(_02835_),
    .A2(_02836_),
    .B(_02262_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08380_ (.I(_02837_),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08381_ (.A1(_00708_),
    .A2(_01378_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08382_ (.I(_02839_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08383_ (.I(_01672_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08384_ (.A1(_01519_),
    .A2(_02841_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08385_ (.A1(_01425_),
    .A2(_02842_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08386_ (.A1(_02262_),
    .A2(_02840_),
    .A3(_02843_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08387_ (.I(_02844_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08388_ (.I(_02845_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08389_ (.I(_02236_),
    .Z(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08390_ (.A1(_02149_),
    .A2(_02211_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _08391_ (.A1(_02159_),
    .A2(_02847_),
    .A3(_02848_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08392_ (.A1(_01396_),
    .A2(_02173_),
    .A3(_02833_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08393_ (.A1(_00750_),
    .A2(_00730_),
    .A3(_02850_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08394_ (.I(_02851_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08395_ (.A1(_02263_),
    .A2(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08396_ (.I(_02853_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08397_ (.A1(_02838_),
    .A2(_02846_),
    .A3(_02849_),
    .A4(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08398_ (.I(_01445_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08399_ (.A1(_01233_),
    .A2(_01360_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08400_ (.A1(_00753_),
    .A2(_02856_),
    .A3(_02857_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08401_ (.I(_00665_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08402_ (.A1(_02859_),
    .A2(_01251_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08403_ (.A1(_02147_),
    .A2(_01403_),
    .A3(_02860_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08404_ (.A1(_01458_),
    .A2(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08405_ (.A1(_02856_),
    .A2(_02862_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08406_ (.A1(_01370_),
    .A2(_01458_),
    .A3(_01400_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08407_ (.A1(_02856_),
    .A2(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08408_ (.A1(_02858_),
    .A2(_02863_),
    .A3(_02865_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08409_ (.A1(_01360_),
    .A2(_02148_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08410_ (.A1(_01402_),
    .A2(_01672_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08411_ (.I(_01422_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08412_ (.A1(_01373_),
    .A2(_01475_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08413_ (.A1(_01412_),
    .A2(_01416_),
    .A3(_01392_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _08414_ (.A1(_02869_),
    .A2(_02870_),
    .A3(_02871_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08415_ (.A1(_02213_),
    .A2(_01411_),
    .A3(_01408_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _08416_ (.A1(_02869_),
    .A2(_02873_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _08417_ (.A1(_01426_),
    .A2(_01427_),
    .A3(_02872_),
    .A4(_02874_),
    .Z(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08418_ (.A1(_02856_),
    .A2(_02867_),
    .A3(_02868_),
    .A4(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08419_ (.I(_00750_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08420_ (.A1(_02877_),
    .A2(_01380_),
    .A3(_01386_),
    .A4(_02873_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08421_ (.A1(_02878_),
    .A2(_02235_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08422_ (.I(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08423_ (.I(_02880_),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08424_ (.A1(_01420_),
    .A2(_02850_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08425_ (.I(_02882_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08426_ (.A1(_02847_),
    .A2(_02883_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08427_ (.A1(_02866_),
    .A2(_02876_),
    .A3(_02881_),
    .A4(_02884_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08428_ (.A1(_02827_),
    .A2(_02855_),
    .A3(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _08429_ (.A1(_01490_),
    .A2(_02822_),
    .A3(_02886_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08430_ (.A1(_02818_),
    .A2(_02887_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08431_ (.I(_02888_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08432_ (.I(_02863_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08433_ (.I(_02890_),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08434_ (.I0(net1),
    .I1(net9),
    .I2(net25),
    .I3(net17),
    .S0(_01436_),
    .S1(_01438_),
    .Z(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08435_ (.I(_00743_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08436_ (.A1(net38),
    .A2(_02893_),
    .B(_00765_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08437_ (.I(_02894_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08438_ (.I(_02865_),
    .Z(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08439_ (.I(_02858_),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08440_ (.I(_02897_),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08441_ (.I(_02865_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08442_ (.I(_02897_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08443_ (.I(_02876_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08444_ (.A1(_00774_),
    .A2(_01382_),
    .B(_00775_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08445_ (.A1(_02902_),
    .A2(_02828_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08446_ (.A1(_02829_),
    .A2(_01554_),
    .A3(_01560_),
    .B(_02903_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08447_ (.A1(_01330_),
    .A2(_01387_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08448_ (.A1(_01388_),
    .A2(_01554_),
    .A3(_01560_),
    .B(_02905_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08449_ (.A1(_02904_),
    .A2(_02906_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08450_ (.I(_02907_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08451_ (.A1(\as2650.debug_psl[0] ),
    .A2(\as2650.debug_psl[3] ),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08452_ (.A1(_02908_),
    .A2(_02909_),
    .B(_02839_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08453_ (.A1(_02908_),
    .A2(_02909_),
    .B(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08454_ (.A1(_01470_),
    .A2(_01810_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08455_ (.A1(_02908_),
    .A2(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08456_ (.A1(_02908_),
    .A2(_02912_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08457_ (.A1(_01456_),
    .A2(_01407_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08458_ (.A1(_02915_),
    .A2(_01378_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08459_ (.A1(_02913_),
    .A2(_02914_),
    .A3(_02916_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08460_ (.A1(_02904_),
    .A2(_02906_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08461_ (.A1(_02214_),
    .A2(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08462_ (.A1(_02904_),
    .A2(_02906_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08463_ (.A1(_01475_),
    .A2(_02918_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08464_ (.A1(_01456_),
    .A2(_02920_),
    .A3(_02921_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08465_ (.A1(_01371_),
    .A2(_01481_),
    .A3(_01377_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08466_ (.A1(_01419_),
    .A2(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08467_ (.I(_02924_),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08468_ (.A1(_02919_),
    .A2(_02922_),
    .B1(_02925_),
    .B2(_02904_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08469_ (.A1(_02911_),
    .A2(_02917_),
    .A3(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08470_ (.I(_02927_),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08471_ (.A1(_02263_),
    .A2(_02835_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08472_ (.I(_02929_),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _08473_ (.A1(_02236_),
    .A2(_02878_),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08474_ (.I(_02931_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08475_ (.A1(_02190_),
    .A2(_02880_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08476_ (.A1(_02187_),
    .A2(_02932_),
    .B(_02933_),
    .C(_02838_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08477_ (.A1(_01332_),
    .A2(_02930_),
    .B(_02934_),
    .C(_02854_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08478_ (.I(_01027_),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08479_ (.A1(_02229_),
    .A2(_02870_),
    .A3(_01524_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08480_ (.A1(_02236_),
    .A2(_02937_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08481_ (.I(_02938_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08482_ (.A1(_02936_),
    .A2(_02939_),
    .B(_02884_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08483_ (.I(_00808_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08484_ (.A1(_01810_),
    .A2(_02941_),
    .B(_02912_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08485_ (.I(_02884_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08486_ (.I(_02876_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08487_ (.A1(_02935_),
    .A2(_02940_),
    .B1(_02942_),
    .B2(_02943_),
    .C(_02944_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08488_ (.A1(_02901_),
    .A2(_02928_),
    .B(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(_02900_),
    .A2(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08490_ (.A1(_01262_),
    .A2(_02898_),
    .B(_02899_),
    .C(_02947_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08491_ (.I(_02863_),
    .Z(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08492_ (.A1(_02895_),
    .A2(_02896_),
    .B(_02948_),
    .C(_02949_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08493_ (.A1(_02891_),
    .A2(_02892_),
    .B(_02950_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08494_ (.I(_02951_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08495_ (.I(_02952_),
    .Z(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08496_ (.I(_02821_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08497_ (.A1(_01426_),
    .A2(_01428_),
    .A3(_02872_),
    .A4(_02874_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08498_ (.I(_02955_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08499_ (.I(_02857_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _08500_ (.I(_02957_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08501_ (.A1(_01365_),
    .A2(_01573_),
    .A3(_02956_),
    .A4(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08502_ (.A1(_02954_),
    .A2(_02959_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08503_ (.I(_01490_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08504_ (.A1(_02961_),
    .A2(_02817_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08505_ (.A1(_02960_),
    .A2(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08506_ (.I(_01366_),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08507_ (.A1(_02818_),
    .A2(_02887_),
    .B(_02963_),
    .C(_02964_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08508_ (.I(_02965_),
    .Z(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08509_ (.I(_02928_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08510_ (.I(_02963_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08511_ (.A1(\as2650.regs[7][0] ),
    .A2(_02966_),
    .B1(_02967_),
    .B2(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08512_ (.A1(_02889_),
    .A2(_02953_),
    .B(_02969_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08513_ (.I0(net2),
    .I1(net10),
    .I2(net26),
    .I3(net18),
    .S0(_01436_),
    .S1(_01438_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08514_ (.A1(_00783_),
    .A2(net131),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08515_ (.A1(net39),
    .A2(net131),
    .B(_02971_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08516_ (.I(_02972_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08517_ (.A1(_00708_),
    .A2(_02173_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08518_ (.A1(_00783_),
    .A2(_01433_),
    .B(_00784_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08519_ (.A1(_02975_),
    .A2(_02830_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08520_ (.I(_02976_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08521_ (.A1(_02936_),
    .A2(_01627_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08522_ (.A1(_01575_),
    .A2(_01576_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08523_ (.A1(_01593_),
    .A2(_01264_),
    .B(_02979_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08524_ (.I(_02829_),
    .Z(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08525_ (.A1(_02978_),
    .A2(_02980_),
    .B(_02981_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08526_ (.A1(_02274_),
    .A2(_02981_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08527_ (.A1(_02978_),
    .A2(_02980_),
    .B(_01389_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _08528_ (.A1(_02977_),
    .A2(_02982_),
    .B1(_02983_),
    .B2(_02984_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08529_ (.I(_01388_),
    .Z(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08530_ (.A1(_01340_),
    .A2(_02986_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08531_ (.A1(_01578_),
    .A2(_02976_),
    .A3(_02987_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08532_ (.A1(_02831_),
    .A2(_01561_),
    .B(_02903_),
    .C(_02906_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08533_ (.A1(_02985_),
    .A2(_02988_),
    .B1(_02989_),
    .B2(_02914_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08534_ (.A1(_02985_),
    .A2(_02988_),
    .Z(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08535_ (.A1(_02914_),
    .A2(_02991_),
    .A3(_02989_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08536_ (.A1(_01574_),
    .A2(_01577_),
    .B(_02986_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08537_ (.A1(_02976_),
    .A2(_02993_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08538_ (.A1(_02907_),
    .A2(_02909_),
    .B(_02918_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08539_ (.A1(_02991_),
    .A2(_02995_),
    .Z(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08540_ (.A1(_02915_),
    .A2(_02173_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08541_ (.A1(_01474_),
    .A2(_02985_),
    .B(_02988_),
    .C(_01372_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08542_ (.A1(_01378_),
    .A2(_02985_),
    .B(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08543_ (.A1(_02924_),
    .A2(_02994_),
    .B1(_02996_),
    .B2(_02997_),
    .C(_02999_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08544_ (.A1(_02974_),
    .A2(_02990_),
    .A3(_02992_),
    .B(_03000_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08545_ (.I(_03001_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08546_ (.A1(_02901_),
    .A2(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08547_ (.A1(_01420_),
    .A2(_02850_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08548_ (.A1(_02264_),
    .A2(_03004_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08549_ (.I(_03005_),
    .Z(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08550_ (.I(_02845_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08551_ (.A1(_01569_),
    .A2(_02880_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08552_ (.A1(_02189_),
    .A2(_02881_),
    .B(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08553_ (.I(_02837_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08554_ (.A1(_01341_),
    .A2(_02930_),
    .B1(_03009_),
    .B2(_03010_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08555_ (.A1(_01483_),
    .A2(_01568_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08556_ (.A1(_02846_),
    .A2(_03012_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08557_ (.A1(_03007_),
    .A2(_03011_),
    .B(_03013_),
    .C(_02939_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08558_ (.I(_02854_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08559_ (.A1(_01588_),
    .A2(_03015_),
    .B(_03006_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08560_ (.I(_01680_),
    .Z(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08561_ (.I(_03017_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08562_ (.I(_03018_),
    .Z(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08563_ (.A1(_01673_),
    .A2(_03019_),
    .A3(_02955_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08564_ (.A1(_02187_),
    .A2(_03006_),
    .B1(_03014_),
    .B2(_03016_),
    .C(_03020_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08565_ (.A1(_03003_),
    .A2(_03021_),
    .B(_02900_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08566_ (.A1(_01264_),
    .A2(_02898_),
    .B(_02865_),
    .C(_03022_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08567_ (.A1(_02973_),
    .A2(_02896_),
    .B(_03023_),
    .C(_02949_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08568_ (.A1(_02891_),
    .A2(_02970_),
    .B(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08569_ (.I(_03025_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08570_ (.I(_03026_),
    .Z(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08571_ (.I(_03002_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08572_ (.A1(\as2650.regs[7][1] ),
    .A2(_02966_),
    .B1(_03028_),
    .B2(_02968_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08573_ (.A1(_02889_),
    .A2(_03027_),
    .B(_03029_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08574_ (.I(\as2650.ext_io_addr[6] ),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08575_ (.I0(net3),
    .I1(net11),
    .I2(net27),
    .I3(net19),
    .S0(_01436_),
    .S1(_03030_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08576_ (.I(_02897_),
    .Z(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08577_ (.I(_02944_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08578_ (.I0(_01384_),
    .I1(_01596_),
    .S(_01388_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08579_ (.I0(_01594_),
    .I1(_01596_),
    .S(_02829_),
    .Z(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _08580_ (.A1(_03034_),
    .A2(_03035_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08581_ (.A1(_01574_),
    .A2(_01577_),
    .B(_02981_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08582_ (.A1(_02976_),
    .A2(_02993_),
    .B1(_02987_),
    .B2(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08583_ (.A1(_02988_),
    .A2(_02995_),
    .B(_03038_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08584_ (.A1(_03036_),
    .A2(_03039_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08585_ (.A1(_02997_),
    .A2(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08586_ (.I(_03034_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08587_ (.A1(_02987_),
    .A2(_03037_),
    .B(_02994_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08588_ (.A1(_02990_),
    .A2(_03043_),
    .B(_03036_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08589_ (.A1(_02990_),
    .A2(_03036_),
    .A3(_03043_),
    .Z(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08590_ (.A1(_03044_),
    .A2(_03045_),
    .Z(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08591_ (.A1(_03034_),
    .A2(_03035_),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08592_ (.A1(_03034_),
    .A2(_03035_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08593_ (.A1(_01474_),
    .A2(_03047_),
    .B(_03048_),
    .C(_01372_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08594_ (.A1(_02214_),
    .A2(_03047_),
    .B(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08595_ (.A1(_02925_),
    .A2(_03042_),
    .B1(_03046_),
    .B2(_02916_),
    .C(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08596_ (.A1(_03041_),
    .A2(_03051_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08597_ (.I(_03052_),
    .Z(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08598_ (.I(_02943_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08599_ (.I(_01077_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08600_ (.I(_02938_),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08601_ (.I(_02884_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08602_ (.I(_02929_),
    .Z(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08603_ (.I(_01048_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08604_ (.I(_02931_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08605_ (.A1(_03059_),
    .A2(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08606_ (.A1(_02186_),
    .A2(_02881_),
    .B(_02837_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08607_ (.A1(_01349_),
    .A2(_03058_),
    .B1(_03061_),
    .B2(_03062_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08608_ (.I(_02844_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08609_ (.A1(_01483_),
    .A2(_01568_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08610_ (.A1(_03059_),
    .A2(_03065_),
    .Z(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08611_ (.A1(_03064_),
    .A2(_03066_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08612_ (.A1(_02846_),
    .A2(_03063_),
    .B(_03067_),
    .C(_02939_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08613_ (.A1(_03055_),
    .A2(_03056_),
    .B(_03057_),
    .C(_03068_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08614_ (.I(_02944_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08615_ (.A1(_01569_),
    .A2(_03054_),
    .B(_03069_),
    .C(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08616_ (.A1(_03033_),
    .A2(_03053_),
    .B(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08617_ (.A1(_01590_),
    .A2(_01055_),
    .B(_01591_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08618_ (.A1(_03073_),
    .A2(_02900_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08619_ (.A1(_02153_),
    .A2(_01374_),
    .A3(_01376_),
    .A4(_01399_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08620_ (.A1(_01365_),
    .A2(_03075_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08621_ (.I(_03076_),
    .Z(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08622_ (.A1(_03032_),
    .A2(_03072_),
    .B(_03074_),
    .C(_03077_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08623_ (.I(_01384_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08624_ (.I(_03079_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08625_ (.I(_03080_),
    .Z(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08626_ (.A1(_03081_),
    .A2(_02896_),
    .B(_02949_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08627_ (.A1(_02891_),
    .A2(_03031_),
    .B1(_03078_),
    .B2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08628_ (.I(_03083_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08629_ (.I(_03084_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08630_ (.I(_03053_),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08631_ (.A1(\as2650.regs[7][2] ),
    .A2(_02966_),
    .B1(_03086_),
    .B2(_02968_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08632_ (.A1(_02889_),
    .A2(_03085_),
    .B(_03087_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08633_ (.I(\as2650.ext_io_addr[7] ),
    .Z(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08634_ (.I0(net4),
    .I1(net12),
    .I2(net28),
    .I3(net20),
    .S0(_03088_),
    .S1(_03030_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08635_ (.I0(net41),
    .I1(net53),
    .S(_01382_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08636_ (.A1(_03090_),
    .A2(_02830_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08637_ (.A1(_02830_),
    .A2(_01606_),
    .B(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08638_ (.A1(_01355_),
    .A2(_02986_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08639_ (.A1(_01389_),
    .A2(_01606_),
    .B(_03093_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08640_ (.A1(_03092_),
    .A2(_03094_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08641_ (.I(_03095_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08642_ (.A1(_03036_),
    .A2(_03039_),
    .B(_03047_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08643_ (.A1(_03096_),
    .A2(_03097_),
    .B(_02839_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08644_ (.A1(_03096_),
    .A2(_03097_),
    .B(_03098_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08645_ (.A1(_03042_),
    .A2(_03035_),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08646_ (.A1(_03044_),
    .A2(_03096_),
    .A3(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08647_ (.A1(_03044_),
    .A2(_03100_),
    .B(_03096_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08648_ (.A1(_02974_),
    .A2(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08649_ (.A1(_03101_),
    .A2(_03103_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08650_ (.I(_03092_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08651_ (.A1(_02925_),
    .A2(_03105_),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08652_ (.I(_03094_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08653_ (.A1(_03105_),
    .A2(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08654_ (.A1(_03105_),
    .A2(_03107_),
    .B(_01372_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08655_ (.A1(_02214_),
    .A2(_03108_),
    .B(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08656_ (.A1(_01476_),
    .A2(_03108_),
    .B(_03110_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08657_ (.A1(_03099_),
    .A2(_03104_),
    .A3(_03106_),
    .A4(_03111_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08658_ (.I(_03112_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08659_ (.A1(_02936_),
    .A2(_03059_),
    .B(_01483_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08660_ (.A1(_01602_),
    .A2(_03114_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08661_ (.A1(_01357_),
    .A2(_02930_),
    .B(_03064_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08662_ (.A1(_03055_),
    .A2(_02932_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08663_ (.A1(_02180_),
    .A2(_03060_),
    .B(_03117_),
    .C(_03010_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08664_ (.A1(_03007_),
    .A2(_03115_),
    .B1(_03116_),
    .B2(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08665_ (.A1(_01613_),
    .A2(_03015_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08666_ (.A1(_03015_),
    .A2(_03119_),
    .B(_03120_),
    .C(_03057_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08667_ (.A1(_01588_),
    .A2(_03054_),
    .B(_03121_),
    .C(_03070_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08668_ (.A1(_03033_),
    .A2(_03113_),
    .B(_03122_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08669_ (.A1(_01074_),
    .A2(_01079_),
    .A3(_02900_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08670_ (.A1(_03032_),
    .A2(_03123_),
    .B(_03124_),
    .C(_03077_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08671_ (.A1(net41),
    .A2(_02893_),
    .B(_00734_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08672_ (.I(_03126_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08673_ (.I(_03127_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08674_ (.A1(_03128_),
    .A2(_02896_),
    .B(_02949_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08675_ (.A1(_02891_),
    .A2(_03089_),
    .B1(_03125_),
    .B2(_03129_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08676_ (.I(_03130_),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08677_ (.I(_03131_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08678_ (.I(_03113_),
    .Z(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08679_ (.A1(\as2650.regs[7][3] ),
    .A2(_02966_),
    .B1(_03133_),
    .B2(_02968_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08680_ (.A1(_02889_),
    .A2(_03132_),
    .B(_03134_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08681_ (.I(_02888_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08682_ (.I(_02863_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08683_ (.I0(net5),
    .I1(net13),
    .I2(net29),
    .I3(net21),
    .S0(_03088_),
    .S1(\as2650.ext_io_addr[6] ),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08684_ (.I(_02172_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08685_ (.I0(_01612_),
    .I1(_02182_),
    .S(_02879_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08686_ (.A1(net207),
    .A2(_03058_),
    .B1(_03139_),
    .B2(_03010_),
    .C(_02853_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08687_ (.A1(_03138_),
    .A2(_02854_),
    .B(_03140_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(_01603_),
    .A2(_03005_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08689_ (.A1(_03006_),
    .A2(_03141_),
    .B(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08690_ (.A1(_00710_),
    .A2(_01433_),
    .B(_00714_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08691_ (.A1(_03144_),
    .A2(_02981_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08692_ (.A1(_02831_),
    .A2(_01618_),
    .B(_03145_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08693_ (.A1(_00658_),
    .A2(_02986_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08694_ (.A1(_01389_),
    .A2(_01618_),
    .B(_03147_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08695_ (.A1(_03146_),
    .A2(_03148_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08696_ (.I(_03149_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08697_ (.A1(_03092_),
    .A2(_03107_),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08698_ (.A1(_03095_),
    .A2(_03097_),
    .B(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08699_ (.A1(_03150_),
    .A2(_03152_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08700_ (.I(_03105_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08701_ (.A1(_03154_),
    .A2(_03107_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08702_ (.A1(_03102_),
    .A2(_03150_),
    .A3(_03155_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08703_ (.A1(_03102_),
    .A2(_03155_),
    .B(_03150_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08704_ (.A1(_02916_),
    .A2(_03156_),
    .A3(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08705_ (.I(_02924_),
    .Z(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08706_ (.I(_03146_),
    .Z(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08707_ (.A1(_03160_),
    .A2(_03148_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08708_ (.A1(_01475_),
    .A2(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08709_ (.A1(_03160_),
    .A2(_03148_),
    .B(_01373_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08710_ (.A1(_01379_),
    .A2(_03161_),
    .B(_03162_),
    .C(_03163_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08711_ (.A1(_03159_),
    .A2(_03160_),
    .B(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _08712_ (.A1(_02840_),
    .A2(_03153_),
    .B(_03158_),
    .C(_03165_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08713_ (.I(_03166_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08714_ (.A1(_02876_),
    .A2(_03167_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08715_ (.A1(_02944_),
    .A2(_03143_),
    .B(_03168_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08716_ (.I0(_01614_),
    .I1(_03169_),
    .S(_02897_),
    .Z(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08717_ (.A1(net42),
    .A2(_02893_),
    .B(_00744_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08718_ (.I(_03171_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08719_ (.A1(_03172_),
    .A2(_03076_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08720_ (.A1(_03076_),
    .A2(_03170_),
    .B(_03173_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08721_ (.A1(_02890_),
    .A2(_03174_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08722_ (.A1(_03136_),
    .A2(_03137_),
    .B(_03175_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08723_ (.I(_03176_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08724_ (.I(_03177_),
    .Z(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08725_ (.I(_02965_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08726_ (.I(_03167_),
    .Z(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08727_ (.I(_02963_),
    .Z(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08728_ (.A1(\as2650.regs[7][4] ),
    .A2(_03179_),
    .B1(_03180_),
    .B2(_03181_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08729_ (.A1(_03135_),
    .A2(_03178_),
    .B(_03182_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08730_ (.I0(net6),
    .I1(net14),
    .I2(net30),
    .I3(net22),
    .S0(\as2650.ext_io_addr[7] ),
    .S1(\as2650.ext_io_addr[6] ),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08731_ (.I(_02925_),
    .Z(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08732_ (.A1(_00717_),
    .A2(_01433_),
    .B(_00718_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08733_ (.A1(_02831_),
    .A2(_01635_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08734_ (.A1(_03185_),
    .A2(_02832_),
    .B(_03186_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08735_ (.A1(_01390_),
    .A2(_01635_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08736_ (.A1(_00650_),
    .A2(_01390_),
    .B(_03188_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08737_ (.A1(_03187_),
    .A2(_03189_),
    .Z(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08738_ (.I(_03160_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08739_ (.A1(_03191_),
    .A2(_03148_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08740_ (.A1(_03157_),
    .A2(_03190_),
    .A3(_03192_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08741_ (.A1(_03157_),
    .A2(_03192_),
    .B(_03190_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08742_ (.A1(_02974_),
    .A2(_03194_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08743_ (.A1(_03193_),
    .A2(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08744_ (.I(_02997_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08745_ (.A1(_03149_),
    .A2(_03152_),
    .B(_03161_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08746_ (.A1(_03190_),
    .A2(_03198_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08747_ (.A1(_03187_),
    .A2(_03189_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08748_ (.A1(_03187_),
    .A2(_03189_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08749_ (.A1(_01411_),
    .A2(_03200_),
    .B(_03201_),
    .C(_01373_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08750_ (.A1(_01481_),
    .A2(_03200_),
    .B(_03202_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08751_ (.A1(_03197_),
    .A2(_03199_),
    .B(_03203_),
    .C(_03159_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08752_ (.A1(_03184_),
    .A2(_03187_),
    .B1(_03196_),
    .B2(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08753_ (.I(_03205_),
    .Z(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08754_ (.I(_00929_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08755_ (.I(_03207_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08756_ (.I(_01626_),
    .Z(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08757_ (.A1(_02177_),
    .A2(_02931_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08758_ (.A1(_03209_),
    .A2(_02932_),
    .B(_03210_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08759_ (.A1(net208),
    .A2(_03058_),
    .B1(_03211_),
    .B2(_03010_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08760_ (.A1(_02226_),
    .A2(_02172_),
    .Z(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08761_ (.A1(_02845_),
    .A2(_03213_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08762_ (.A1(_03064_),
    .A2(_03212_),
    .B(_03214_),
    .C(_02938_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08763_ (.A1(_03208_),
    .A2(_03056_),
    .B(_02943_),
    .C(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08764_ (.A1(_01613_),
    .A2(_03057_),
    .B(_03216_),
    .C(_02901_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08765_ (.A1(_03070_),
    .A2(_03206_),
    .B(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08766_ (.A1(_00753_),
    .A2(_01446_),
    .A3(_02957_),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08767_ (.A1(_01630_),
    .A2(_03219_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08768_ (.A1(_02898_),
    .A2(_03218_),
    .B(_03220_),
    .C(_03077_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08769_ (.A1(_00717_),
    .A2(_01434_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08770_ (.A1(net34),
    .A2(_01434_),
    .B(_03222_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08771_ (.I(_03223_),
    .Z(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08772_ (.A1(_03224_),
    .A2(_02899_),
    .B(_02890_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _08773_ (.A1(_03136_),
    .A2(_03183_),
    .B1(_03221_),
    .B2(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08774_ (.I(_03226_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08775_ (.I(_03227_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08776_ (.I(_03206_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08777_ (.A1(\as2650.regs[7][5] ),
    .A2(_03179_),
    .B1(_03229_),
    .B2(_03181_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08778_ (.A1(_03135_),
    .A2(_03228_),
    .B(_03230_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08779_ (.I0(net7),
    .I1(net15),
    .I2(net31),
    .I3(net23),
    .S0(_03088_),
    .S1(_03030_),
    .Z(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08780_ (.A1(_00701_),
    .A2(_01434_),
    .B(_00706_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08781_ (.A1(_02832_),
    .A2(_01647_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08782_ (.A1(_03232_),
    .A2(_02832_),
    .B(_03233_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08783_ (.I(_02916_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08784_ (.A1(_01390_),
    .A2(_01648_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08785_ (.A1(_00642_),
    .A2(_01391_),
    .B(_03236_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08786_ (.A1(_03234_),
    .A2(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08787_ (.A1(_03234_),
    .A2(_03237_),
    .Z(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08788_ (.A1(_03238_),
    .A2(_03239_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08789_ (.A1(_03185_),
    .A2(_02833_),
    .B(_03186_),
    .C(_03189_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08790_ (.A1(_03194_),
    .A2(_03240_),
    .A3(_03241_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08791_ (.A1(_03194_),
    .A2(_03241_),
    .B(_03240_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08792_ (.A1(_03235_),
    .A2(_03242_),
    .A3(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08793_ (.A1(_03200_),
    .A2(_03198_),
    .B(_03201_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08794_ (.A1(_03240_),
    .A2(_03245_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08795_ (.A1(_01481_),
    .A2(_03239_),
    .B1(_03240_),
    .B2(_01379_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08796_ (.A1(_03197_),
    .A2(_03246_),
    .B1(_03247_),
    .B2(_01374_),
    .C(_03159_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08797_ (.A1(_03184_),
    .A2(_03234_),
    .B1(_03244_),
    .B2(_03248_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08798_ (.I(_03249_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08799_ (.I(_02941_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(_02171_),
    .A2(_02880_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08801_ (.A1(_03208_),
    .A2(_02932_),
    .B(_02837_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08802_ (.A1(net209),
    .A2(_03058_),
    .B1(_03252_),
    .B2(_03253_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08803_ (.A1(_02226_),
    .A2(_02172_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08804_ (.A1(_03207_),
    .A2(_03255_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08805_ (.A1(_02845_),
    .A2(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08806_ (.A1(_02846_),
    .A2(_03254_),
    .B(_03257_),
    .C(_02938_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08807_ (.A1(_03251_),
    .A2(_03056_),
    .B(_02943_),
    .C(_03258_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08808_ (.A1(_03138_),
    .A2(_03054_),
    .B(_03259_),
    .C(_02901_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08809_ (.A1(_03033_),
    .A2(_03250_),
    .B(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08810_ (.A1(_00990_),
    .A2(_03219_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08811_ (.A1(_03032_),
    .A2(_03261_),
    .B(_03262_),
    .C(_03077_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08812_ (.A1(net35),
    .A2(_02893_),
    .B(_00727_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08813_ (.I(_03264_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08814_ (.I(_03265_),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08815_ (.A1(_03266_),
    .A2(_02899_),
    .B(_02890_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08816_ (.A1(_03136_),
    .A2(_03231_),
    .B1(_03263_),
    .B2(_03267_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08817_ (.I(_03268_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08818_ (.I(_03269_),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08819_ (.I(_03250_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08820_ (.A1(\as2650.regs[7][6] ),
    .A2(_03179_),
    .B1(_03271_),
    .B2(_03181_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08821_ (.A1(_03135_),
    .A2(_03270_),
    .B(_03272_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _08822_ (.I0(net8),
    .I1(net16),
    .I2(net32),
    .I3(net24),
    .S0(_03088_),
    .S1(_03030_),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08823_ (.A1(_00723_),
    .A2(net131),
    .B(_00724_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08824_ (.I(_03274_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08825_ (.A1(_03275_),
    .A2(_02864_),
    .B(_02862_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08826_ (.A1(_01367_),
    .A2(_03276_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08827_ (.I0(_01677_),
    .I1(_01657_),
    .S(_01391_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08828_ (.I0(_01653_),
    .I1(_01657_),
    .S(_02833_),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08829_ (.A1(_03278_),
    .A2(_03279_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08830_ (.A1(_03278_),
    .A2(_03279_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08831_ (.A1(_03280_),
    .A2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08832_ (.I(_03237_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08833_ (.A1(_03234_),
    .A2(_03283_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08834_ (.A1(_03243_),
    .A2(_03282_),
    .A3(_03284_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08835_ (.A1(_03243_),
    .A2(_03284_),
    .B(_03282_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08836_ (.A1(_02974_),
    .A2(_03285_),
    .A3(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08837_ (.I(_03238_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08838_ (.A1(_03288_),
    .A2(_03245_),
    .B(_03239_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08839_ (.A1(_03282_),
    .A2(_03289_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08840_ (.A1(_02840_),
    .A2(_03290_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08841_ (.A1(_01476_),
    .A2(_03281_),
    .B1(_03282_),
    .B2(_02160_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08842_ (.I(_03159_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _08843_ (.A1(_01457_),
    .A2(_03292_),
    .B(_03293_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08844_ (.A1(_03287_),
    .A2(_03291_),
    .A3(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08845_ (.A1(_03184_),
    .A2(_03278_),
    .B(_03295_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08846_ (.I(_03296_),
    .Z(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08847_ (.I(_01810_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08848_ (.I(_01057_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08849_ (.A1(_03298_),
    .A2(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08850_ (.A1(_02912_),
    .A2(_03300_),
    .Z(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08851_ (.A1(_03251_),
    .A2(_03060_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08852_ (.A1(_02166_),
    .A2(_02881_),
    .B(_02838_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08853_ (.A1(net210),
    .A2(_02930_),
    .B1(_03302_),
    .B2(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08854_ (.A1(_03207_),
    .A2(_03209_),
    .B(_02226_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08855_ (.A1(_02941_),
    .A2(_03305_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08856_ (.A1(_03064_),
    .A2(_03306_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _08857_ (.A1(_03007_),
    .A2(_03304_),
    .B(_03307_),
    .C(_02939_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08858_ (.A1(_03056_),
    .A2(_03301_),
    .B(_03308_),
    .C(_03057_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08859_ (.A1(_01642_),
    .A2(_03054_),
    .B(_03309_),
    .C(_03070_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08860_ (.A1(_03033_),
    .A2(_03297_),
    .B(_03310_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08861_ (.A1(_01654_),
    .A2(_02898_),
    .B(_02899_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08862_ (.A1(_03032_),
    .A2(_03311_),
    .B(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08863_ (.A1(_03136_),
    .A2(_03273_),
    .B1(_03277_),
    .B2(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08864_ (.I(_03314_),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08865_ (.I(_03315_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08866_ (.I(_03297_),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08867_ (.A1(\as2650.regs[7][7] ),
    .A2(_03179_),
    .B1(_03317_),
    .B2(_03181_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08868_ (.A1(_03135_),
    .A2(_03316_),
    .B(_03318_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08869_ (.A1(_02592_),
    .A2(_02480_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08870_ (.I(_03319_),
    .Z(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08871_ (.I0(_02548_),
    .I1(\as2650.stack[1][0] ),
    .S(_03320_),
    .Z(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08872_ (.I(_03321_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08873_ (.I0(_02553_),
    .I1(\as2650.stack[1][1] ),
    .S(_03320_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08874_ (.I(_03322_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08875_ (.I0(_02555_),
    .I1(\as2650.stack[1][2] ),
    .S(_03320_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08876_ (.I(_03323_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08877_ (.I0(_02557_),
    .I1(\as2650.stack[1][3] ),
    .S(_03320_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08878_ (.I(_03324_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08879_ (.I(_03319_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08880_ (.I0(_02559_),
    .I1(\as2650.stack[1][4] ),
    .S(_03325_),
    .Z(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08881_ (.I(_03326_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08882_ (.I0(_02562_),
    .I1(\as2650.stack[1][5] ),
    .S(_03325_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08883_ (.I(_03327_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08884_ (.I0(_02564_),
    .I1(\as2650.stack[1][6] ),
    .S(_03325_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08885_ (.I(_03328_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08886_ (.I0(_02566_),
    .I1(\as2650.stack[1][7] ),
    .S(_03325_),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08887_ (.I(_03329_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08888_ (.I(_03319_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08889_ (.I0(_02568_),
    .I1(\as2650.stack[1][8] ),
    .S(_03330_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08890_ (.I(_03331_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08891_ (.I0(_02571_),
    .I1(\as2650.stack[1][9] ),
    .S(_03330_),
    .Z(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08892_ (.I(_03332_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08893_ (.I0(_02573_),
    .I1(\as2650.stack[1][10] ),
    .S(_03330_),
    .Z(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08894_ (.I(_03333_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08895_ (.I0(_02575_),
    .I1(\as2650.stack[1][11] ),
    .S(_03330_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08896_ (.I(_03334_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08897_ (.I(_03319_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08898_ (.I0(_02577_),
    .I1(\as2650.stack[1][12] ),
    .S(_03335_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08899_ (.I(_03336_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08900_ (.I0(_02580_),
    .I1(\as2650.stack[1][13] ),
    .S(_03335_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08901_ (.I(_03337_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08902_ (.I0(_02582_),
    .I1(\as2650.stack[1][14] ),
    .S(_03335_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08903_ (.I(_03338_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08904_ (.I0(_02584_),
    .I1(\as2650.stack[1][15] ),
    .S(_03335_),
    .Z(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08905_ (.I(_03339_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08906_ (.I(_01551_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08907_ (.A1(\as2650.last_addr[0] ),
    .A2(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08908_ (.A1(_01566_),
    .A2(_03341_),
    .B(_01692_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08909_ (.A1(_01287_),
    .A2(net214),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08910_ (.A1(\as2650.last_addr[1] ),
    .A2(_01552_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08911_ (.A1(_01450_),
    .A2(_03342_),
    .A3(_03343_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08912_ (.I(_01691_),
    .Z(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08913_ (.A1(\as2650.last_addr[2] ),
    .A2(_01589_),
    .B(_01599_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08914_ (.A1(_03344_),
    .A2(_03345_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08915_ (.A1(_01295_),
    .A2(net214),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08916_ (.A1(\as2650.last_addr[3] ),
    .A2(_03340_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08917_ (.A1(_01450_),
    .A2(_03346_),
    .A3(_03347_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_01303_),
    .A2(_01583_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08919_ (.A1(\as2650.last_addr[4] ),
    .A2(_01571_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08920_ (.A1(_03348_),
    .A2(_03349_),
    .B(_01692_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08921_ (.A1(\as2650.last_addr[5] ),
    .A2(_03340_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08922_ (.A1(_01450_),
    .A2(_01640_),
    .A3(_03350_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08923_ (.A1(_01316_),
    .A2(_01583_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(\as2650.last_addr[6] ),
    .A2(_01571_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08925_ (.A1(_03351_),
    .A2(_03352_),
    .B(_01692_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08926_ (.I(_01462_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08927_ (.A1(\as2650.last_addr[7] ),
    .A2(_03340_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08928_ (.A1(_03353_),
    .A2(_01662_),
    .A3(_03354_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08929_ (.I(_01542_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08930_ (.I(\as2650.indirect_target[0] ),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08931_ (.I(_01362_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08932_ (.I(_03356_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08933_ (.I(_01368_),
    .Z(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08934_ (.I(_03358_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08935_ (.I(_01424_),
    .Z(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08936_ (.I(_01683_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08937_ (.A1(_02144_),
    .A2(_03360_),
    .A3(_03361_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08938_ (.I(_03362_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08939_ (.I(_03363_),
    .Z(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08940_ (.I(_02902_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08941_ (.I(_03365_),
    .Z(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08942_ (.I(_00747_),
    .Z(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08943_ (.I(_01522_),
    .Z(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08944_ (.A1(_02205_),
    .A2(_03367_),
    .A3(_03368_),
    .A4(_01668_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08945_ (.A1(_03360_),
    .A2(_03361_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08946_ (.A1(_01671_),
    .A2(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08947_ (.I(_02206_),
    .Z(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08948_ (.A1(_03372_),
    .A2(_03371_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08949_ (.A1(_01686_),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08950_ (.I(_03374_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08951_ (.I(_00957_),
    .Z(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08952_ (.A1(_01359_),
    .A2(_01363_),
    .A3(_02148_),
    .B(\as2650.instruction_args_latch[8] ),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08953_ (.A1(_03365_),
    .A2(_01664_),
    .A3(_01444_),
    .A4(_01404_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08954_ (.A1(_03377_),
    .A2(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08955_ (.A1(_03376_),
    .A2(_03379_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08956_ (.A1(_03366_),
    .A2(_03369_),
    .A3(_03371_),
    .B1(_03375_),
    .B2(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08957_ (.A1(_01675_),
    .A2(_01684_),
    .A3(_02823_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08958_ (.I(_03382_),
    .Z(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08959_ (.A1(_01676_),
    .A2(_03381_),
    .B1(_03383_),
    .B2(_03355_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08960_ (.I(_02825_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08961_ (.A1(_03385_),
    .A2(_03370_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08962_ (.I(\as2650.instruction_args_latch[0] ),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08963_ (.I(_00960_),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08964_ (.A1(_03388_),
    .A2(_01663_),
    .A3(_01444_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08965_ (.I(_03389_),
    .Z(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08966_ (.I(_03390_),
    .Z(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08967_ (.I(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08968_ (.A1(_02143_),
    .A2(_02902_),
    .A3(_01358_),
    .A4(_01363_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08969_ (.A1(_03387_),
    .A2(_03392_),
    .B(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08970_ (.A1(_03364_),
    .A2(_03384_),
    .B1(_03386_),
    .B2(_03394_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08971_ (.A1(_03355_),
    .A2(_03357_),
    .B(_03359_),
    .C(_03395_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08972_ (.I(\as2650.indirect_target[1] ),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08973_ (.I(_03382_),
    .Z(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08974_ (.A1(_02213_),
    .A2(_03361_),
    .A3(_01684_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08975_ (.A1(_03377_),
    .A2(_03378_),
    .B(_02223_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _08976_ (.A1(_01359_),
    .A2(_01364_),
    .A3(_02148_),
    .B(\as2650.instruction_args_latch[9] ),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08977_ (.I(_02975_),
    .Z(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08978_ (.A1(_03401_),
    .A2(_01664_),
    .A3(_01445_),
    .A4(_01405_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08979_ (.A1(_03400_),
    .A2(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08980_ (.I(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _08981_ (.A1(_02287_),
    .A2(_03399_),
    .A3(_03404_),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08982_ (.I(_02206_),
    .Z(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08983_ (.A1(_03372_),
    .A2(_03405_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08984_ (.A1(_02972_),
    .A2(_03406_),
    .B(_03407_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08985_ (.I(_03371_),
    .Z(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08986_ (.A1(_03398_),
    .A2(_03405_),
    .B1(_03408_),
    .B2(_03409_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08987_ (.A1(_03396_),
    .A2(_03397_),
    .B1(_03410_),
    .B2(_01676_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08988_ (.A1(_02144_),
    .A2(_01358_),
    .A3(_01363_),
    .B(\as2650.instruction_args_latch[1] ),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08989_ (.A1(_03388_),
    .A2(_03401_),
    .A3(_01664_),
    .A4(_01444_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08990_ (.A1(_03412_),
    .A2(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08991_ (.I(_03386_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08992_ (.A1(_03364_),
    .A2(_03411_),
    .B1(_03414_),
    .B2(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08993_ (.A1(_03396_),
    .A2(_03357_),
    .B(_03359_),
    .C(_03416_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08994_ (.I(\as2650.indirect_target[2] ),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08995_ (.I(\as2650.instruction_args_latch[10] ),
    .Z(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08996_ (.I0(_00738_),
    .I1(_03418_),
    .S(_01679_),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08997_ (.I(_03419_),
    .Z(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08998_ (.A1(_02287_),
    .A2(_03400_),
    .A3(_03402_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08999_ (.A1(_03400_),
    .A2(_03402_),
    .B(_02287_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09000_ (.A1(_03399_),
    .A2(_03421_),
    .B(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09001_ (.A1(_02300_),
    .A2(_03420_),
    .A3(_03423_),
    .Z(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09002_ (.A1(_03372_),
    .A2(_03424_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09003_ (.A1(_03080_),
    .A2(_03406_),
    .B(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09004_ (.A1(_03398_),
    .A2(_03424_),
    .B1(_03426_),
    .B2(_03409_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09005_ (.A1(_03417_),
    .A2(_03397_),
    .B1(_03427_),
    .B2(_01676_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09006_ (.I0(_00738_),
    .I1(\as2650.instruction_args_latch[2] ),
    .S(_03389_),
    .Z(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09007_ (.A1(_03364_),
    .A2(_03428_),
    .B1(_03429_),
    .B2(_03415_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09008_ (.A1(_03417_),
    .A2(_03357_),
    .B(_03359_),
    .C(_03430_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09009_ (.I(\as2650.indirect_target[3] ),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09010_ (.A1(\as2650.instruction_args_latch[11] ),
    .A2(_01680_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09011_ (.A1(_03126_),
    .A2(_03017_),
    .B(_03432_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09012_ (.A1(_02297_),
    .A2(_02299_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09013_ (.A1(_03434_),
    .A2(_03419_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09014_ (.A1(_03434_),
    .A2(_03420_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09015_ (.A1(_03435_),
    .A2(_03423_),
    .B(_03436_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09016_ (.A1(_02308_),
    .A2(_03433_),
    .A3(_03437_),
    .Z(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09017_ (.I(_02206_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09018_ (.I(_03439_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09019_ (.I(_03372_),
    .Z(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09020_ (.A1(_03441_),
    .A2(_03438_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09021_ (.A1(_03128_),
    .A2(_03440_),
    .B(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09022_ (.I(_03371_),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09023_ (.A1(_03398_),
    .A2(_03438_),
    .B1(_03443_),
    .B2(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09024_ (.I(_01675_),
    .Z(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09025_ (.I(_03446_),
    .Z(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09026_ (.A1(_03431_),
    .A2(_03397_),
    .B1(_03445_),
    .B2(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(\as2650.instruction_args_latch[3] ),
    .A2(_03389_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09028_ (.A1(_03126_),
    .A2(_03389_),
    .B(_03449_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09029_ (.I(_03386_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09030_ (.A1(_03364_),
    .A2(_03448_),
    .B1(_03450_),
    .B2(_03451_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09031_ (.A1(_03431_),
    .A2(_03357_),
    .B(_03359_),
    .C(_03452_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09032_ (.I(\as2650.indirect_target[4] ),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09033_ (.I(_03356_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09034_ (.I(_03358_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09035_ (.I(_03362_),
    .Z(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09036_ (.I(_03144_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09037_ (.I(_01680_),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09038_ (.A1(\as2650.instruction_args_latch[12] ),
    .A2(_03458_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09039_ (.A1(_03171_),
    .A2(_03458_),
    .B(_03459_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09040_ (.I(_03460_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09041_ (.A1(_02308_),
    .A2(_03433_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09042_ (.A1(_02308_),
    .A2(_03433_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09043_ (.A1(_03462_),
    .A2(_03437_),
    .B(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09044_ (.A1(_02326_),
    .A2(_03461_),
    .A3(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09045_ (.A1(_03457_),
    .A2(_03369_),
    .A3(_03444_),
    .B1(_03375_),
    .B2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09046_ (.A1(_03453_),
    .A2(_03397_),
    .B1(_03466_),
    .B2(_03447_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09047_ (.A1(\as2650.instruction_args_latch[4] ),
    .A2(_03390_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09048_ (.A1(_03171_),
    .A2(_03391_),
    .B(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09049_ (.A1(_03456_),
    .A2(_03467_),
    .B1(_03469_),
    .B2(_03451_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09050_ (.A1(_03453_),
    .A2(_03454_),
    .B(_03455_),
    .C(_03470_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09051_ (.I(\as2650.indirect_target[5] ),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09052_ (.I(_03382_),
    .Z(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(_00748_),
    .A2(_03458_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09054_ (.A1(_03223_),
    .A2(_03018_),
    .B(_03473_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09055_ (.A1(_02324_),
    .A2(_03460_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09056_ (.A1(_02325_),
    .A2(_03460_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09057_ (.A1(_03475_),
    .A2(_03464_),
    .B(_03476_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09058_ (.A1(_02341_),
    .A2(_03474_),
    .A3(_03477_),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09059_ (.A1(_03439_),
    .A2(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09060_ (.A1(_03224_),
    .A2(_03441_),
    .B(_03479_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09061_ (.A1(_03398_),
    .A2(_03478_),
    .B1(_03480_),
    .B2(_03444_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09062_ (.A1(_03471_),
    .A2(_03472_),
    .B1(_03481_),
    .B2(_03447_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09063_ (.A1(\as2650.instruction_args_latch[5] ),
    .A2(_03390_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09064_ (.A1(_03223_),
    .A2(_03391_),
    .B(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09065_ (.A1(_03456_),
    .A2(_03482_),
    .B1(_03484_),
    .B2(_03451_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09066_ (.A1(_03471_),
    .A2(_03454_),
    .B(_03455_),
    .C(_03485_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09067_ (.I(\as2650.indirect_target[6] ),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09068_ (.A1(_03266_),
    .A2(_03439_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09069_ (.I(_03487_),
    .Z(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09070_ (.I(_03232_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09071_ (.A1(_00756_),
    .A2(_03017_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09072_ (.A1(_03489_),
    .A2(_03017_),
    .B(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09073_ (.A1(_02356_),
    .A2(_03491_),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09074_ (.A1(_02341_),
    .A2(_03474_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09075_ (.A1(_02340_),
    .A2(_03474_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09076_ (.A1(_03493_),
    .A2(_03477_),
    .B(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09077_ (.A1(_03492_),
    .A2(_03495_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09078_ (.A1(_03409_),
    .A2(_03488_),
    .B1(_03496_),
    .B2(_03375_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09079_ (.A1(_03486_),
    .A2(_03472_),
    .B1(_03497_),
    .B2(_03447_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09080_ (.A1(\as2650.instruction_args_latch[6] ),
    .A2(_03392_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09081_ (.A1(_03264_),
    .A2(_03392_),
    .B(_03499_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09082_ (.A1(_03456_),
    .A2(_03498_),
    .B1(_03500_),
    .B2(_03451_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09083_ (.A1(_03486_),
    .A2(_03454_),
    .B(_03455_),
    .C(_03501_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09084_ (.I(\as2650.indirect_target[7] ),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09085_ (.I(net315),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09086_ (.A1(\as2650.instruction_args_latch[14] ),
    .A2(_03458_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09087_ (.A1(_03264_),
    .A2(_03018_),
    .B(_03504_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09088_ (.I(_03505_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09089_ (.A1(_02356_),
    .A2(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09090_ (.I(_03492_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09091_ (.A1(_03493_),
    .A2(_03477_),
    .B(_03508_),
    .C(_03494_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09092_ (.A1(_03507_),
    .A2(_03509_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09093_ (.A1(_02369_),
    .A2(_03503_),
    .A3(_03510_),
    .Z(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09094_ (.A1(_03409_),
    .A2(_03488_),
    .B1(_03511_),
    .B2(_03375_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09095_ (.A1(_03502_),
    .A2(_03472_),
    .B1(_03512_),
    .B2(_03446_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09096_ (.A1(\as2650.instruction_args_latch[7] ),
    .A2(_03391_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09097_ (.A1(_01678_),
    .A2(_03392_),
    .B(_03514_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09098_ (.A1(_03456_),
    .A2(_03513_),
    .B1(_03515_),
    .B2(_03386_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09099_ (.A1(_03502_),
    .A2(_03454_),
    .B(_03455_),
    .C(_03516_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09100_ (.I(\as2650.indirect_target[8] ),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09101_ (.I(_01367_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09102_ (.I(_03518_),
    .Z(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09103_ (.I(_03519_),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09104_ (.A1(_02383_),
    .A2(_03506_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09105_ (.A1(_02383_),
    .A2(_03505_),
    .Z(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09106_ (.A1(_03521_),
    .A2(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09107_ (.A1(_02381_),
    .A2(_02368_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09108_ (.A1(_03524_),
    .A2(_03506_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(_03524_),
    .A2(_03506_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09110_ (.A1(_03509_),
    .A2(_03525_),
    .B(_03526_),
    .C(_03507_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09111_ (.A1(_03523_),
    .A2(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09112_ (.A1(_03444_),
    .A2(_03488_),
    .B1(_03528_),
    .B2(_03374_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09113_ (.A1(_03517_),
    .A2(_03472_),
    .B1(_03529_),
    .B2(_03446_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09114_ (.A1(_03379_),
    .A2(_03415_),
    .B1(_03530_),
    .B2(_03363_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09115_ (.A1(_03517_),
    .A2(_01455_),
    .B(_03520_),
    .C(_03531_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09116_ (.I(_01362_),
    .Z(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09117_ (.I(_03532_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09118_ (.A1(_03388_),
    .A2(_01665_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09119_ (.A1(_03360_),
    .A2(_03361_),
    .A3(_03534_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09120_ (.I(_03535_),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09121_ (.A1(_02398_),
    .A2(_03491_),
    .Z(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09122_ (.I(_03505_),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09123_ (.A1(_02383_),
    .A2(_03538_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09124_ (.A1(_03522_),
    .A2(_03527_),
    .B(_03539_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09125_ (.A1(_03537_),
    .A2(_03540_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09126_ (.I(_03374_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09127_ (.A1(_03446_),
    .A2(_03542_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09128_ (.I(_03382_),
    .Z(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09129_ (.A1(\as2650.indirect_target[9] ),
    .A2(_03544_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09130_ (.A1(_03541_),
    .A2(_03543_),
    .B(_03545_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09131_ (.I(_03388_),
    .Z(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09132_ (.I(_03370_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09133_ (.A1(_03547_),
    .A2(_03548_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09134_ (.A1(\as2650.indirect_target[9] ),
    .A2(_03533_),
    .B1(_03536_),
    .B2(_03403_),
    .C1(_03546_),
    .C2(_03549_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09135_ (.A1(_03344_),
    .A2(_03550_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09136_ (.I(_03535_),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09137_ (.A1(_02412_),
    .A2(_03491_),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09138_ (.A1(_03523_),
    .A2(_03537_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09139_ (.A1(_02399_),
    .A2(_03538_),
    .B1(_03527_),
    .B2(_03553_),
    .C(_03539_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09140_ (.A1(_03552_),
    .A2(_03554_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09141_ (.A1(\as2650.indirect_target[10] ),
    .A2(_03544_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09142_ (.A1(_03543_),
    .A2(_03555_),
    .B(_03556_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09143_ (.A1(\as2650.indirect_target[10] ),
    .A2(_03533_),
    .B1(_03551_),
    .B2(_03420_),
    .C1(_03557_),
    .C2(_03549_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09144_ (.A1(_03344_),
    .A2(_03558_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09145_ (.I(_01460_),
    .Z(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09146_ (.I(_03433_),
    .Z(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09147_ (.I(_01666_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09148_ (.A1(_03561_),
    .A2(_01674_),
    .A3(_03374_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09149_ (.I(_03562_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09150_ (.A1(_02426_),
    .A2(_03503_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09151_ (.A1(_02413_),
    .A2(_03538_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09152_ (.I(_03538_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09153_ (.A1(_02413_),
    .A2(_03566_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09154_ (.A1(_03565_),
    .A2(_03554_),
    .B(_03567_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09155_ (.A1(_03564_),
    .A2(_03568_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09156_ (.A1(\as2650.indirect_target[11] ),
    .A2(_03544_),
    .B1(_03563_),
    .B2(_03569_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09157_ (.A1(_03363_),
    .A2(_03570_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09158_ (.A1(\as2650.indirect_target[11] ),
    .A2(_03533_),
    .B1(_03536_),
    .B2(_03560_),
    .C(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09159_ (.A1(_03559_),
    .A2(_03572_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_02413_),
    .A2(_02426_),
    .B(_03566_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09161_ (.A1(_03552_),
    .A2(_03554_),
    .A3(_03564_),
    .B(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09162_ (.A1(_02439_),
    .A2(_03566_),
    .A3(_03574_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09163_ (.A1(\as2650.indirect_target[12] ),
    .A2(_03544_),
    .B1(_03562_),
    .B2(_03575_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09164_ (.A1(_03363_),
    .A2(_03576_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09165_ (.A1(\as2650.indirect_target[12] ),
    .A2(_03533_),
    .B1(_03536_),
    .B2(_03461_),
    .C(_03577_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09166_ (.A1(_03559_),
    .A2(_03578_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09167_ (.I(_01446_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09168_ (.I(_03579_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09169_ (.I(_03535_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09170_ (.A1(\as2650.indirect_target[13] ),
    .A2(_03383_),
    .B1(_03563_),
    .B2(_02446_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09171_ (.I(_03367_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09172_ (.I(_03185_),
    .Z(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09173_ (.I(_03584_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09174_ (.A1(_00760_),
    .A2(_03019_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09175_ (.A1(_03585_),
    .A2(_03019_),
    .B(_03586_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09176_ (.A1(_03367_),
    .A2(_03587_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09177_ (.A1(_02446_),
    .A2(_03583_),
    .B(_03551_),
    .C(_03588_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09178_ (.A1(_03581_),
    .A2(_03582_),
    .B(_03589_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09179_ (.A1(_03580_),
    .A2(_03590_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09180_ (.I(_03591_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09181_ (.A1(\as2650.indirect_target[14] ),
    .A2(_03383_),
    .B1(_03563_),
    .B2(_02454_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09182_ (.A1(_03367_),
    .A2(_03503_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09183_ (.A1(_02454_),
    .A2(_03583_),
    .B(_03551_),
    .C(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09184_ (.A1(_03536_),
    .A2(_03592_),
    .B(_03594_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09185_ (.A1(_03580_),
    .A2(_03595_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09186_ (.I(_03596_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09187_ (.A1(_03581_),
    .A2(_03563_),
    .B(_02462_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09188_ (.A1(\as2650.indirect_target[15] ),
    .A2(_03383_),
    .A3(_03415_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09189_ (.I(_01691_),
    .Z(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09190_ (.A1(_03597_),
    .A2(_03598_),
    .B(_03599_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09191_ (.I(_00925_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09192_ (.I(_00739_),
    .Z(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09193_ (.A1(_03601_),
    .A2(_03551_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09194_ (.A1(_03600_),
    .A2(_03581_),
    .B1(_03602_),
    .B2(\as2650.indexed_cyc[0] ),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09195_ (.A1(_03579_),
    .A2(_02958_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09196_ (.I(_03604_),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09197_ (.A1(_03603_),
    .A2(_03605_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09198_ (.I(_00759_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09199_ (.A1(_03606_),
    .A2(_03581_),
    .B1(_03602_),
    .B2(\as2650.indexed_cyc[1] ),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09200_ (.A1(_03605_),
    .A2(_03607_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09201_ (.I(_01405_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09202_ (.A1(_03360_),
    .A2(_01674_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09203_ (.A1(_00677_),
    .A2(_03547_),
    .B1(_03608_),
    .B2(_03609_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09204_ (.A1(_03532_),
    .A2(_03610_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09205_ (.A1(_01170_),
    .A2(_01381_),
    .B1(_03548_),
    .B2(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09206_ (.A1(_03605_),
    .A2(_03612_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09207_ (.I(_03519_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09208_ (.I(_01533_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09209_ (.I(_03614_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09210_ (.I(_03615_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09211_ (.I(_03616_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09212_ (.I(_02230_),
    .Z(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09213_ (.A1(_03618_),
    .A2(_02870_),
    .A3(_02871_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09214_ (.A1(_03617_),
    .A2(_03619_),
    .B(net205),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09215_ (.I(_01665_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09216_ (.A1(_01276_),
    .A2(_03621_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09217_ (.A1(_03613_),
    .A2(_03620_),
    .A3(_03622_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09218_ (.A1(_01193_),
    .A2(_02146_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09219_ (.I(_02868_),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09220_ (.A1(_03624_),
    .A2(_02151_),
    .B(_03608_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09221_ (.A1(_03623_),
    .A2(_03625_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09222_ (.I(_03615_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09223_ (.I(_02836_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09224_ (.A1(_02869_),
    .A2(_01457_),
    .A3(_02841_),
    .A4(_02158_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09225_ (.A1(_03628_),
    .A2(_03629_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09226_ (.A1(_01422_),
    .A2(_02213_),
    .A3(_02841_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _09227_ (.A1(_02205_),
    .A2(_02160_),
    .A3(_01521_),
    .A4(_03631_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09228_ (.A1(_02869_),
    .A2(_02201_),
    .A3(_01393_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09229_ (.A1(_03197_),
    .A2(_03631_),
    .B(_03632_),
    .C(_03633_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09230_ (.A1(_03630_),
    .A2(_03634_),
    .B(_01669_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09231_ (.I(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09232_ (.I(_03636_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09233_ (.A1(_03627_),
    .A2(_03637_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09234_ (.A1(_03632_),
    .A2(_03638_),
    .B(_01462_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09235_ (.A1(_03621_),
    .A2(_03626_),
    .B1(_03638_),
    .B2(_02877_),
    .C(_03639_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09236_ (.I(\as2650.warmup[1] ),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09237_ (.A1(\as2650.warmup[0] ),
    .A2(_03640_),
    .B(_01260_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09238_ (.A1(\as2650.warmup[0] ),
    .A2(\as2650.warmup[1] ),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09239_ (.A1(_01260_),
    .A2(_03641_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09240_ (.I(_03385_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09241_ (.I(_03642_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09242_ (.I(_03385_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09243_ (.A1(_03601_),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09244_ (.I(_03645_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09245_ (.A1(_03366_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(\as2650.instruction_args_latch[0] ),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09246_ (.A1(_03605_),
    .A2(_03647_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09247_ (.I(_03604_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09248_ (.I(_03648_),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09249_ (.I(_03401_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09250_ (.A1(_03650_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(\as2650.instruction_args_latch[1] ),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09251_ (.A1(_03649_),
    .A2(_03651_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09252_ (.I(_00738_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09253_ (.I(_03652_),
    .Z(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09254_ (.A1(_03653_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(\as2650.instruction_args_latch[2] ),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09255_ (.A1(_03649_),
    .A2(_03654_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09256_ (.I(_03090_),
    .Z(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09257_ (.A1(_03655_),
    .A2(_03643_),
    .B1(_03646_),
    .B2(\as2650.instruction_args_latch[3] ),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09258_ (.A1(_03649_),
    .A2(_03656_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09259_ (.I(_03644_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09260_ (.I(_03645_),
    .Z(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09261_ (.A1(_03457_),
    .A2(_03657_),
    .B1(_03658_),
    .B2(\as2650.instruction_args_latch[4] ),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09262_ (.A1(_03649_),
    .A2(_03659_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09263_ (.I(_03585_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09264_ (.A1(_03660_),
    .A2(_03657_),
    .B1(_03658_),
    .B2(\as2650.instruction_args_latch[5] ),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09265_ (.A1(_03648_),
    .A2(_03661_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09266_ (.I(_03489_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09267_ (.A1(_03662_),
    .A2(_03657_),
    .B1(_03658_),
    .B2(\as2650.instruction_args_latch[6] ),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09268_ (.A1(_03648_),
    .A2(_03663_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09269_ (.A1(_03275_),
    .A2(_03657_),
    .B1(_03658_),
    .B2(\as2650.instruction_args_latch[7] ),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09270_ (.A1(_03648_),
    .A2(_03664_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09271_ (.I(_02957_),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09272_ (.I(_02867_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09273_ (.A1(_03666_),
    .A2(_03622_),
    .Z(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09274_ (.A1(_03601_),
    .A2(_03665_),
    .A3(_03667_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09275_ (.I(_03668_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09276_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09277_ (.I(_03667_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(_03366_),
    .A2(_03671_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09279_ (.A1(_03670_),
    .A2(_03672_),
    .B(_03599_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09280_ (.A1(\as2650.instruction_args_latch[9] ),
    .A2(_03669_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09281_ (.A1(_03650_),
    .A2(_03671_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09282_ (.A1(_03673_),
    .A2(_03674_),
    .B(_03599_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09283_ (.A1(_03653_),
    .A2(_03671_),
    .B1(_03669_),
    .B2(_03418_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09284_ (.A1(_03559_),
    .A2(_03675_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09285_ (.A1(_03655_),
    .A2(_03671_),
    .B1(_03669_),
    .B2(\as2650.instruction_args_latch[11] ),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09286_ (.A1(_03559_),
    .A2(_03676_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09287_ (.I(_01691_),
    .Z(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09288_ (.I(_03667_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09289_ (.I(_03668_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09290_ (.A1(_03457_),
    .A2(_03678_),
    .B1(_03679_),
    .B2(\as2650.instruction_args_latch[12] ),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09291_ (.A1(_03677_),
    .A2(_03680_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09292_ (.A1(_03660_),
    .A2(_03678_),
    .B1(_03679_),
    .B2(_00748_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09293_ (.A1(_03677_),
    .A2(_03681_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09294_ (.A1(_03662_),
    .A2(_03678_),
    .B1(_03679_),
    .B2(\as2650.instruction_args_latch[14] ),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09295_ (.A1(_03677_),
    .A2(_03682_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09296_ (.A1(_03275_),
    .A2(_03678_),
    .B1(_03679_),
    .B2(\as2650.instruction_args_latch[15] ),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09297_ (.A1(_03677_),
    .A2(_03683_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09298_ (.I(_02153_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09299_ (.A1(_01674_),
    .A2(_02150_),
    .B(_03608_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09300_ (.I(_02848_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09301_ (.I(_03686_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09302_ (.I(_03687_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09303_ (.A1(_02872_),
    .A2(_03635_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09304_ (.A1(_03688_),
    .A2(_03689_),
    .B(_03601_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09305_ (.A1(_03623_),
    .A2(_03685_),
    .A3(_03690_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09306_ (.A1(_03684_),
    .A2(_03627_),
    .A3(_03642_),
    .B1(_03691_),
    .B2(_03532_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09307_ (.I(_02860_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09308_ (.A1(_01370_),
    .A2(_01376_),
    .B(_03693_),
    .C(_03622_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09309_ (.A1(_01376_),
    .A2(_03692_),
    .B(_03694_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09310_ (.A1(net48),
    .A2(net47),
    .A3(net49),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09311_ (.A1(net44),
    .A2(net43),
    .A3(net46),
    .A4(net45),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09312_ (.A1(_01375_),
    .A2(_00672_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09313_ (.A1(_00739_),
    .A2(_01361_),
    .B1(_03698_),
    .B2(_02859_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09314_ (.A1(_03696_),
    .A2(_03697_),
    .B(_01897_),
    .C(_03699_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09315_ (.I(_03700_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09316_ (.A1(_03684_),
    .A2(_03693_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09317_ (.A1(_01361_),
    .A2(_02155_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09318_ (.I(_03703_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09319_ (.A1(_03358_),
    .A2(_03704_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09320_ (.A1(_03695_),
    .A2(_03701_),
    .A3(_03702_),
    .A4(_03705_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09321_ (.I(_03706_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09322_ (.I(_01403_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09323_ (.I(_03534_),
    .Z(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09324_ (.I(_02234_),
    .Z(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09325_ (.I(_03709_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09326_ (.I(_03710_),
    .Z(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09327_ (.A1(_03561_),
    .A2(_01670_),
    .B1(_02872_),
    .B2(_03711_),
    .C(_00664_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(_03625_),
    .A2(_03712_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09329_ (.A1(_03583_),
    .A2(_03708_),
    .A3(_03548_),
    .B1(_03713_),
    .B2(_03547_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09330_ (.A1(_03707_),
    .A2(_03356_),
    .B1(_03693_),
    .B2(_00672_),
    .C1(_03714_),
    .C2(_01233_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09331_ (.A1(_03579_),
    .A2(_02861_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09332_ (.A1(_02153_),
    .A2(_03707_),
    .A3(_02859_),
    .A4(_01251_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09333_ (.I(_03717_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09334_ (.A1(_03716_),
    .A2(_03718_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09335_ (.A1(_01185_),
    .A2(_01455_),
    .B(_03701_),
    .C(_03719_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09336_ (.A1(_03715_),
    .A2(_03720_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09337_ (.A1(_01375_),
    .A2(_03532_),
    .B(_03707_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09338_ (.A1(_01399_),
    .A2(_03619_),
    .B(_01251_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09339_ (.A1(_03707_),
    .A2(_03722_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09340_ (.A1(_03621_),
    .A2(_03723_),
    .B(_02859_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09341_ (.A1(_00676_),
    .A2(_03721_),
    .B1(_03724_),
    .B2(_03684_),
    .C(_03701_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09342_ (.A1(_01463_),
    .A2(_03725_),
    .Z(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09343_ (.I(_03726_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09344_ (.I(_02842_),
    .Z(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09345_ (.A1(_02197_),
    .A2(_03631_),
    .A3(_03235_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09346_ (.A1(_01428_),
    .A2(_02867_),
    .A3(_03624_),
    .A4(_03728_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09347_ (.A1(_01476_),
    .A2(_01523_),
    .A3(_03727_),
    .A4(_03729_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09348_ (.I(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09349_ (.A1(_03684_),
    .A2(_02154_),
    .A3(_03621_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09350_ (.I(_03732_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09351_ (.A1(_01375_),
    .A2(_03731_),
    .B(_03733_),
    .C(_02861_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09352_ (.A1(_03622_),
    .A2(_03700_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09353_ (.A1(_03734_),
    .A2(_03735_),
    .B(_03599_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09354_ (.I(_02895_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09355_ (.I(_01529_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09356_ (.I(_03737_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09357_ (.I(_03738_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09358_ (.I(_03739_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09359_ (.I(_03740_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09360_ (.A1(\as2650.insin[0] ),
    .A2(_03617_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09361_ (.I(_03519_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09362_ (.A1(_03736_),
    .A2(_03741_),
    .B(_03742_),
    .C(_03743_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09363_ (.I(_02973_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09364_ (.A1(\as2650.insin[1] ),
    .A2(_03617_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09365_ (.A1(_03744_),
    .A2(_03741_),
    .B(_03745_),
    .C(_03743_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09366_ (.A1(\as2650.insin[2] ),
    .A2(_03617_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09367_ (.I(_03518_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09368_ (.I(_03747_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09369_ (.A1(_03081_),
    .A2(_03741_),
    .B(_03746_),
    .C(_03748_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09370_ (.I(_03128_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09371_ (.I(_03616_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09372_ (.A1(\as2650.insin[3] ),
    .A2(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09373_ (.A1(_03749_),
    .A2(_03741_),
    .B(_03751_),
    .C(_03748_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09374_ (.I(_03172_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09375_ (.I(_03752_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09376_ (.I(_03740_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09377_ (.A1(\as2650.insin[4] ),
    .A2(_03750_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09378_ (.A1(_03753_),
    .A2(_03754_),
    .B(_03755_),
    .C(_03748_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09379_ (.I(_03224_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09380_ (.A1(\as2650.insin[5] ),
    .A2(_03750_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09381_ (.A1(_03756_),
    .A2(_03754_),
    .B(_03757_),
    .C(_03748_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _09382_ (.I(_03266_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09383_ (.A1(\as2650.insin[6] ),
    .A2(_03750_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09384_ (.I(_03747_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09385_ (.A1(_03758_),
    .A2(_03754_),
    .B(_03759_),
    .C(_03760_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09386_ (.I(_01678_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09387_ (.I(_03761_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09388_ (.A1(\as2650.insin[7] ),
    .A2(_03740_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09389_ (.A1(_03762_),
    .A2(_03754_),
    .B(_03763_),
    .C(_03760_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09390_ (.I(_03703_),
    .Z(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09391_ (.I(_03764_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09392_ (.I(_03765_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09393_ (.A1(_02145_),
    .A2(_02212_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09394_ (.I(_03767_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09395_ (.A1(_02825_),
    .A2(_03768_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09396_ (.I(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09397_ (.I(_03770_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09398_ (.I(_01533_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09399_ (.A1(_02209_),
    .A2(_03727_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09400_ (.I(_03773_),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09401_ (.A1(_03772_),
    .A2(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09402_ (.I(_03775_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09403_ (.A1(\as2650.debug_psu[3] ),
    .A2(_02526_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09404_ (.I(_03777_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09405_ (.I(_03778_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09406_ (.I(_03779_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09407_ (.I(_03780_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09408_ (.I(_03781_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09409_ (.A1(\as2650.debug_psu[0] ),
    .A2(_01861_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09410_ (.A1(_02247_),
    .A2(_03783_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09411_ (.I(_03784_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09412_ (.I(_03785_),
    .Z(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09413_ (.I(_03786_),
    .Z(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09414_ (.I(_02258_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09415_ (.I(_03783_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09416_ (.I(_03789_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09417_ (.I(_03790_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09418_ (.I(_03791_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09419_ (.I(_03792_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09420_ (.A1(\as2650.stack[2][13] ),
    .A2(_03788_),
    .B1(_03793_),
    .B2(\as2650.stack[3][13] ),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09421_ (.I(_02474_),
    .Z(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09422_ (.I(_02590_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09423_ (.A1(\as2650.stack[1][13] ),
    .A2(_03795_),
    .B1(_03796_),
    .B2(\as2650.stack[0][13] ),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09424_ (.A1(_03787_),
    .A2(_03794_),
    .A3(_03797_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09425_ (.A1(_01868_),
    .A2(_03783_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09426_ (.I(_03799_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09427_ (.I(_03800_),
    .Z(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09428_ (.I(_03801_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09429_ (.I(_03802_),
    .Z(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09430_ (.I(_02474_),
    .Z(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09431_ (.I(_02590_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09432_ (.A1(\as2650.stack[5][13] ),
    .A2(_03804_),
    .B1(_03805_),
    .B2(\as2650.stack[4][13] ),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09433_ (.I(_03792_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09434_ (.A1(\as2650.stack[6][13] ),
    .A2(_03788_),
    .B1(_03807_),
    .B2(\as2650.stack[7][13] ),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09435_ (.A1(_03803_),
    .A2(_03806_),
    .A3(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09436_ (.A1(_03782_),
    .A2(_03798_),
    .A3(_03809_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09437_ (.I(_03777_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09438_ (.I(_03811_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09439_ (.I(_03812_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09440_ (.I(_03787_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09441_ (.A1(\as2650.stack[10][13] ),
    .A2(_03788_),
    .B1(_03793_),
    .B2(\as2650.stack[11][13] ),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09442_ (.A1(\as2650.stack[9][13] ),
    .A2(_03795_),
    .B1(_03796_),
    .B2(\as2650.stack[8][13] ),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09443_ (.A1(_03814_),
    .A2(_03815_),
    .A3(_03816_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09444_ (.A1(\as2650.stack[13][13] ),
    .A2(_03795_),
    .B1(_03796_),
    .B2(\as2650.stack[12][13] ),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09445_ (.A1(\as2650.stack[14][13] ),
    .A2(_03788_),
    .B1(_03793_),
    .B2(\as2650.stack[15][13] ),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09446_ (.A1(_03803_),
    .A2(_03818_),
    .A3(_03819_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09447_ (.A1(_03813_),
    .A2(_03817_),
    .A3(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09448_ (.A1(_03810_),
    .A2(_03821_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09449_ (.A1(_03609_),
    .A2(_03767_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09450_ (.I(_03823_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09451_ (.A1(_03666_),
    .A2(_03824_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09452_ (.A1(_03369_),
    .A2(_03825_),
    .B(_03776_),
    .C(_02446_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09453_ (.A1(_03776_),
    .A2(_03822_),
    .B(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09454_ (.A1(_03377_),
    .A2(_03378_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09455_ (.A1(_03080_),
    .A2(_03018_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09456_ (.A1(_03418_),
    .A2(_03019_),
    .B(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09457_ (.I(_02203_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09458_ (.I(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09459_ (.A1(net203),
    .A2(_03832_),
    .B(_03500_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09460_ (.A1(net200),
    .A2(_03831_),
    .B(_03469_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09461_ (.A1(net198),
    .A2(_02204_),
    .B(_03429_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09462_ (.A1(net196),
    .A2(_02202_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09463_ (.A1(_03387_),
    .A2(_03390_),
    .B(_03393_),
    .C(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09464_ (.A1(net197),
    .A2(_02203_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09465_ (.A1(_03412_),
    .A2(_03413_),
    .A3(_03838_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09466_ (.A1(_03412_),
    .A2(_03413_),
    .B(_03838_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09467_ (.A1(_03837_),
    .A2(_03839_),
    .B(_03840_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09468_ (.A1(net198),
    .A2(_02204_),
    .A3(_03429_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09469_ (.A1(_03835_),
    .A2(_03841_),
    .B(_03842_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09470_ (.A1(net199),
    .A2(_02203_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09471_ (.A1(_03450_),
    .A2(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09472_ (.A1(net199),
    .A2(_02204_),
    .A3(_03450_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09473_ (.A1(_03843_),
    .A2(_03845_),
    .B(_03846_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09474_ (.A1(net200),
    .A2(_03832_),
    .A3(_03469_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09475_ (.A1(_03834_),
    .A2(_03847_),
    .B(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09476_ (.A1(net201),
    .A2(_03831_),
    .A3(_03484_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09477_ (.A1(net201),
    .A2(_03831_),
    .B(_03484_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09478_ (.A1(_03850_),
    .A2(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09479_ (.A1(_03849_),
    .A2(_03852_),
    .B(_03850_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09480_ (.I(_03832_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09481_ (.A1(net203),
    .A2(_03854_),
    .A3(_03500_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09482_ (.A1(_03833_),
    .A2(_03853_),
    .B(_03855_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09483_ (.I(_03515_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(net204),
    .A2(_03832_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09485_ (.A1(_03857_),
    .A2(_03858_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09486_ (.A1(_03857_),
    .A2(_03858_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09487_ (.A1(_03856_),
    .A2(_03859_),
    .B(_03860_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09488_ (.A1(_03828_),
    .A2(_03404_),
    .A3(_03830_),
    .A4(_03861_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09489_ (.A1(_03560_),
    .A2(_03461_),
    .A3(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09490_ (.A1(_03587_),
    .A2(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09491_ (.A1(_03863_),
    .A2(_03587_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09492_ (.A1(_03864_),
    .A2(_03770_),
    .A3(_03865_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09493_ (.I(_03703_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09494_ (.A1(_03771_),
    .A2(_03827_),
    .B(_03866_),
    .C(_03867_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09495_ (.A1(_00760_),
    .A2(_03766_),
    .B(_03868_),
    .C(_03760_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09496_ (.A1(_02823_),
    .A2(_02212_),
    .A3(_03534_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09497_ (.I(_03869_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09498_ (.A1(_03566_),
    .A2(_03864_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09499_ (.I(_02867_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09500_ (.I(_03872_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09501_ (.A1(_03609_),
    .A2(_03768_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09502_ (.I(_03874_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09503_ (.A1(_03441_),
    .A2(_03875_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09504_ (.A1(_02454_),
    .A2(_03873_),
    .A3(_03876_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09505_ (.I(_02258_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09506_ (.A1(\as2650.stack[2][14] ),
    .A2(_03878_),
    .B1(_03807_),
    .B2(\as2650.stack[3][14] ),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09507_ (.A1(\as2650.stack[1][14] ),
    .A2(_03804_),
    .B1(_03805_),
    .B2(\as2650.stack[0][14] ),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09508_ (.A1(_03787_),
    .A2(_03879_),
    .A3(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09509_ (.A1(\as2650.stack[5][14] ),
    .A2(_02474_),
    .B1(_02590_),
    .B2(\as2650.stack[4][14] ),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09510_ (.A1(\as2650.stack[6][14] ),
    .A2(_03878_),
    .B1(_03792_),
    .B2(\as2650.stack[7][14] ),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09511_ (.A1(_03802_),
    .A2(_03882_),
    .A3(_03883_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09512_ (.A1(_03782_),
    .A2(_03881_),
    .A3(_03884_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09513_ (.A1(\as2650.stack[10][14] ),
    .A2(_03878_),
    .B1(_03807_),
    .B2(\as2650.stack[11][14] ),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09514_ (.A1(\as2650.stack[9][14] ),
    .A2(_03804_),
    .B1(_03805_),
    .B2(\as2650.stack[8][14] ),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09515_ (.A1(_03787_),
    .A2(_03886_),
    .A3(_03887_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09516_ (.A1(\as2650.stack[13][14] ),
    .A2(_03804_),
    .B1(_03805_),
    .B2(\as2650.stack[12][14] ),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09517_ (.A1(\as2650.stack[14][14] ),
    .A2(_03878_),
    .B1(_03807_),
    .B2(\as2650.stack[15][14] ),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09518_ (.A1(_03802_),
    .A2(_03889_),
    .A3(_03890_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09519_ (.A1(_03813_),
    .A2(_03888_),
    .A3(_03891_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09520_ (.A1(_03885_),
    .A2(_03892_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09521_ (.A1(\as2650.page_reg[1] ),
    .A2(_03775_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09522_ (.A1(_03776_),
    .A2(_03893_),
    .B(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09523_ (.A1(_03825_),
    .A2(_03895_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09524_ (.I(_03869_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09525_ (.A1(_03877_),
    .A2(_03896_),
    .B(_03897_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09526_ (.A1(_03870_),
    .A2(_03871_),
    .B(_03898_),
    .C(_03867_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09527_ (.A1(_00756_),
    .A2(_03766_),
    .B(_03899_),
    .C(_03760_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09528_ (.A1(_03587_),
    .A2(_03503_),
    .A3(_03863_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09529_ (.I0(_01682_),
    .I1(\as2650.page_reg[2] ),
    .S(_01222_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09530_ (.A1(_03900_),
    .A2(_03901_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09531_ (.I(_03872_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09532_ (.A1(_02462_),
    .A2(_03903_),
    .A3(_03876_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09533_ (.I(_02258_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09534_ (.I(_03792_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09535_ (.A1(\as2650.stack[2][15] ),
    .A2(_03905_),
    .B1(_03906_),
    .B2(\as2650.stack[3][15] ),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09536_ (.A1(\as2650.stack[1][15] ),
    .A2(_02475_),
    .B1(_02591_),
    .B2(\as2650.stack[0][15] ),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09537_ (.A1(_03814_),
    .A2(_03907_),
    .A3(_03908_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09538_ (.A1(\as2650.stack[5][15] ),
    .A2(_03795_),
    .B1(_03796_),
    .B2(\as2650.stack[4][15] ),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09539_ (.A1(\as2650.stack[6][15] ),
    .A2(_03905_),
    .B1(_03793_),
    .B2(\as2650.stack[7][15] ),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09540_ (.A1(_03803_),
    .A2(_03910_),
    .A3(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09541_ (.A1(_03782_),
    .A2(_03909_),
    .A3(_03912_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09542_ (.A1(\as2650.stack[10][15] ),
    .A2(_03905_),
    .B1(_03906_),
    .B2(\as2650.stack[11][15] ),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09543_ (.A1(\as2650.stack[9][15] ),
    .A2(_02475_),
    .B1(_02591_),
    .B2(\as2650.stack[8][15] ),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09544_ (.A1(_03814_),
    .A2(_03914_),
    .A3(_03915_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09545_ (.A1(\as2650.stack[13][15] ),
    .A2(_02475_),
    .B1(_02591_),
    .B2(\as2650.stack[12][15] ),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09546_ (.A1(\as2650.stack[14][15] ),
    .A2(_03905_),
    .B1(_03906_),
    .B2(\as2650.stack[15][15] ),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09547_ (.A1(_03803_),
    .A2(_03917_),
    .A3(_03918_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09548_ (.A1(_03813_),
    .A2(_03916_),
    .A3(_03919_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09549_ (.A1(_03913_),
    .A2(_03920_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(_02462_),
    .A2(_03775_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09551_ (.A1(_03776_),
    .A2(_03921_),
    .B(_03922_),
    .ZN(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09552_ (.A1(_03825_),
    .A2(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09553_ (.I(_03869_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09554_ (.A1(_03904_),
    .A2(_03924_),
    .B(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09555_ (.I(_03764_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09556_ (.A1(_03870_),
    .A2(_03902_),
    .B(_03926_),
    .C(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09557_ (.I(_03732_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09558_ (.I(_01462_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09559_ (.A1(\as2650.instruction_args_latch[15] ),
    .A2(_03929_),
    .B(_03930_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09560_ (.A1(_03928_),
    .A2(_03931_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09561_ (.I(_01254_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09562_ (.A1(\as2650.last_addr[8] ),
    .A2(_03932_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09563_ (.I(_03358_),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09564_ (.A1(_01562_),
    .A2(_03933_),
    .B(_03934_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09565_ (.A1(\as2650.last_addr[9] ),
    .A2(_03932_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09566_ (.A1(_03353_),
    .A2(_01580_),
    .A3(_03935_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09567_ (.A1(\as2650.last_addr[10] ),
    .A2(_03932_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09568_ (.A1(_01597_),
    .A2(_03936_),
    .B(_03934_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09569_ (.A1(\as2650.last_addr[11] ),
    .A2(_03932_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09570_ (.A1(_03353_),
    .A2(_01607_),
    .A3(_03937_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(\as2650.last_addr[12] ),
    .A2(_01643_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09572_ (.A1(_01620_),
    .A2(_03938_),
    .B(_03934_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09573_ (.I(\as2650.last_addr[13] ),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09574_ (.A1(_03939_),
    .A2(net213),
    .B(_03353_),
    .C(_01637_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09575_ (.A1(_01246_),
    .A2(_01643_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(\as2650.last_addr[14] ),
    .A2(_01643_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09577_ (.A1(_03940_),
    .A2(_03941_),
    .B(_03934_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09578_ (.I(\as2650.last_addr[15] ),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09579_ (.A1(_03942_),
    .A2(net213),
    .B(_03580_),
    .C(_01659_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09580_ (.A1(_01519_),
    .A2(_02815_),
    .A3(_02195_),
    .A4(_01526_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09581_ (.A1(_03710_),
    .A2(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09582_ (.I(_03944_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09583_ (.I(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09584_ (.I(_03945_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09585_ (.A1(\as2650.ivectors_base[0] ),
    .A2(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09586_ (.I(_03747_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09587_ (.A1(_02316_),
    .A2(_03946_),
    .B(_03948_),
    .C(_03949_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09588_ (.A1(\as2650.ivectors_base[1] ),
    .A2(_03947_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09589_ (.A1(_02333_),
    .A2(_03946_),
    .B(_03950_),
    .C(_03949_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09590_ (.A1(\as2650.ivectors_base[2] ),
    .A2(_03947_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09591_ (.A1(_02348_),
    .A2(_03946_),
    .B(_03951_),
    .C(_03949_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09592_ (.A1(\as2650.ivectors_base[3] ),
    .A2(_03947_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09593_ (.A1(_02364_),
    .A2(_03946_),
    .B(_03952_),
    .C(_03949_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09594_ (.I(_03945_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09595_ (.I(_03944_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09596_ (.A1(\as2650.ivectors_base[4] ),
    .A2(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09597_ (.I(_03747_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09598_ (.A1(_02375_),
    .A2(_03953_),
    .B(_03955_),
    .C(_03956_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09599_ (.A1(\as2650.ivectors_base[5] ),
    .A2(_03954_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09600_ (.A1(_02393_),
    .A2(_03953_),
    .B(_03957_),
    .C(_03956_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09601_ (.A1(\as2650.ivectors_base[6] ),
    .A2(_03954_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09602_ (.A1(_02406_),
    .A2(_03953_),
    .B(_03958_),
    .C(_03956_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09603_ (.A1(\as2650.ivectors_base[7] ),
    .A2(_03954_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09604_ (.A1(_02421_),
    .A2(_03953_),
    .B(_03959_),
    .C(_03956_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09605_ (.I(_03945_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09606_ (.I(_03944_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09607_ (.A1(\as2650.ivectors_base[8] ),
    .A2(_03961_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09608_ (.I(_03518_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09609_ (.I(_03963_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09610_ (.A1(_02433_),
    .A2(_03960_),
    .B(_03962_),
    .C(_03964_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09611_ (.A1(\as2650.ivectors_base[9] ),
    .A2(_03961_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09612_ (.A1(_02448_),
    .A2(_03960_),
    .B(_03965_),
    .C(_03964_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09613_ (.A1(\as2650.ivectors_base[10] ),
    .A2(_03961_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09614_ (.A1(_02456_),
    .A2(_03960_),
    .B(_03966_),
    .C(_03964_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09615_ (.A1(\as2650.ivectors_base[11] ),
    .A2(_03961_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09616_ (.A1(_02464_),
    .A2(_03960_),
    .B(_03967_),
    .C(_03964_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09617_ (.I(_03708_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09618_ (.I(_01227_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09619_ (.I(_03969_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09620_ (.I(_03768_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09621_ (.A1(_03376_),
    .A2(_03970_),
    .B(_03971_),
    .ZN(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09622_ (.A1(_00681_),
    .A2(_03708_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09623_ (.I(_00953_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09624_ (.I(_03823_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09625_ (.A1(_02895_),
    .A2(_03439_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09626_ (.A1(_03406_),
    .A2(_03380_),
    .B(_03823_),
    .C(_03976_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09627_ (.A1(_02223_),
    .A2(_03974_),
    .A3(_03975_),
    .B(_03977_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09628_ (.A1(_01668_),
    .A2(_03687_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09629_ (.A1(_03376_),
    .A2(_03979_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09630_ (.I(_03773_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09631_ (.I(_03784_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09632_ (.I(_03982_),
    .Z(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09633_ (.I(_02255_),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09634_ (.I(_03984_),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09635_ (.I(_03789_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09636_ (.I(_03986_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09637_ (.A1(\as2650.stack[2][0] ),
    .A2(_03985_),
    .B1(_03987_),
    .B2(\as2650.stack[3][0] ),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09638_ (.I(_02471_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09639_ (.I(_03989_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09640_ (.I(_02587_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09641_ (.I(_03991_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09642_ (.A1(\as2650.stack[1][0] ),
    .A2(_03990_),
    .B1(_03992_),
    .B2(\as2650.stack[0][0] ),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09643_ (.A1(_03983_),
    .A2(_03988_),
    .A3(_03993_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09644_ (.I(_03989_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09645_ (.I(_03991_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09646_ (.A1(\as2650.stack[5][0] ),
    .A2(_03995_),
    .B1(_03996_),
    .B2(\as2650.stack[4][0] ),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09647_ (.I(_03984_),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09648_ (.I(_03986_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09649_ (.A1(\as2650.stack[6][0] ),
    .A2(_03998_),
    .B1(_03999_),
    .B2(\as2650.stack[7][0] ),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09650_ (.A1(_03801_),
    .A2(_03997_),
    .A3(_04000_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09651_ (.A1(_03780_),
    .A2(_03994_),
    .A3(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09652_ (.I(_03811_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09653_ (.A1(\as2650.stack[10][0] ),
    .A2(_03985_),
    .B1(_03987_),
    .B2(\as2650.stack[11][0] ),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09654_ (.A1(\as2650.stack[9][0] ),
    .A2(_03990_),
    .B1(_03992_),
    .B2(\as2650.stack[8][0] ),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09655_ (.A1(_03983_),
    .A2(_04004_),
    .A3(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09656_ (.I(_03799_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09657_ (.I(_04007_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09658_ (.A1(\as2650.stack[13][0] ),
    .A2(_03990_),
    .B1(_03992_),
    .B2(\as2650.stack[12][0] ),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09659_ (.A1(\as2650.stack[14][0] ),
    .A2(_03985_),
    .B1(_03987_),
    .B2(\as2650.stack[15][0] ),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09660_ (.A1(_04008_),
    .A2(_04009_),
    .A3(_04010_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09661_ (.A1(_04003_),
    .A2(_04006_),
    .A3(_04011_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09662_ (.A1(_04002_),
    .A2(_04012_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09663_ (.A1(_03981_),
    .A2(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09664_ (.A1(_03376_),
    .A2(_03774_),
    .B(_04014_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09665_ (.I0(_03980_),
    .I1(_04015_),
    .S(_03637_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09666_ (.I(_03709_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09667_ (.A1(_02223_),
    .A2(_04017_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09668_ (.A1(_03711_),
    .A2(_04016_),
    .B(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09669_ (.I(_01227_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09670_ (.I(_04020_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09671_ (.I(_03872_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09672_ (.A1(_04021_),
    .A2(_03975_),
    .B(_04022_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09673_ (.A1(_03873_),
    .A2(_03978_),
    .B1(_04019_),
    .B2(_04023_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09674_ (.A1(_03968_),
    .A2(_03972_),
    .B1(_03973_),
    .B2(_04024_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09675_ (.A1(_03394_),
    .A2(_03836_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(_03925_),
    .A2(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09677_ (.A1(_04025_),
    .A2(_04027_),
    .B(_03765_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09678_ (.I(_03963_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09679_ (.A1(_03736_),
    .A2(_03766_),
    .B(_04028_),
    .C(_04029_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09680_ (.I(_03764_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09681_ (.A1(_03414_),
    .A2(_03838_),
    .A3(_03837_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09682_ (.I(_03768_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09683_ (.I(_00953_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09684_ (.A1(_04033_),
    .A2(_02288_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09685_ (.A1(_04032_),
    .A2(_04034_),
    .B(_03644_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09686_ (.A1(_00681_),
    .A2(_03534_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09687_ (.I(_03561_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09688_ (.I(_03635_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09689_ (.I(_04038_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09690_ (.I(_02848_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09691_ (.I(_04040_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09692_ (.A1(_00957_),
    .A2(_01423_),
    .A3(_01667_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09693_ (.A1(_02280_),
    .A2(_04042_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09694_ (.A1(_02280_),
    .A2(_04042_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09695_ (.A1(_04043_),
    .A2(_04044_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09696_ (.I(_04040_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09697_ (.A1(_02288_),
    .A2(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09698_ (.A1(_04041_),
    .A2(_04045_),
    .B(_04047_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09699_ (.A1(_02209_),
    .A2(_03727_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09700_ (.I(_04049_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09701_ (.I(_03779_),
    .Z(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09702_ (.I(_03982_),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09703_ (.I(_03984_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09704_ (.I(_03790_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09705_ (.A1(\as2650.stack[2][1] ),
    .A2(_04053_),
    .B1(_04054_),
    .B2(\as2650.stack[3][1] ),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09706_ (.I(_03989_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09707_ (.I(_03991_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09708_ (.A1(\as2650.stack[1][1] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[0][1] ),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09709_ (.A1(_04052_),
    .A2(_04055_),
    .A3(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09710_ (.I(_02472_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09711_ (.I(_02588_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09712_ (.A1(\as2650.stack[5][1] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(\as2650.stack[4][1] ),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09713_ (.I(_02256_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09714_ (.I(_03986_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09715_ (.A1(\as2650.stack[6][1] ),
    .A2(_04063_),
    .B1(_04064_),
    .B2(\as2650.stack[7][1] ),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09716_ (.A1(_04008_),
    .A2(_04062_),
    .A3(_04065_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09717_ (.A1(_04051_),
    .A2(_04059_),
    .A3(_04066_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09718_ (.A1(\as2650.stack[10][1] ),
    .A2(_04063_),
    .B1(_04054_),
    .B2(\as2650.stack[11][1] ),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09719_ (.A1(\as2650.stack[9][1] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(\as2650.stack[8][1] ),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09720_ (.A1(_04052_),
    .A2(_04068_),
    .A3(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09721_ (.I(_04007_),
    .Z(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09722_ (.A1(\as2650.stack[13][1] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(\as2650.stack[12][1] ),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09723_ (.A1(\as2650.stack[14][1] ),
    .A2(_04063_),
    .B1(_04054_),
    .B2(\as2650.stack[15][1] ),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09724_ (.A1(_04071_),
    .A2(_04072_),
    .A3(_04073_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09725_ (.A1(_04003_),
    .A2(_04070_),
    .A3(_04074_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09726_ (.A1(_04067_),
    .A2(_04075_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09727_ (.I(_04049_),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09728_ (.A1(_02288_),
    .A2(_04077_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09729_ (.I(_04038_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09730_ (.A1(_04050_),
    .A2(_04076_),
    .B(_04078_),
    .C(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09731_ (.A1(_04039_),
    .A2(_04048_),
    .B(_04080_),
    .C(_03737_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09732_ (.A1(_02280_),
    .A2(_03614_),
    .B(_04081_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09733_ (.A1(_04037_),
    .A2(_04082_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09734_ (.A1(_03408_),
    .A2(_03824_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09735_ (.I(_04020_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09736_ (.A1(_04085_),
    .A2(_04082_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09737_ (.I(_03874_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09738_ (.A1(_04034_),
    .A2(_04086_),
    .B(_04087_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09739_ (.A1(_03873_),
    .A2(_04084_),
    .A3(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09740_ (.A1(_04036_),
    .A2(_04083_),
    .A3(_04089_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09741_ (.A1(_03897_),
    .A2(_04031_),
    .B1(_04035_),
    .B2(_04090_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09742_ (.A1(_04030_),
    .A2(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09743_ (.A1(_03744_),
    .A2(_03766_),
    .B(_04092_),
    .C(_04029_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09744_ (.I(_03765_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09745_ (.A1(net198),
    .A2(_03854_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09746_ (.A1(_03429_),
    .A2(_04094_),
    .A3(_03841_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09747_ (.A1(_04033_),
    .A2(_02300_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09748_ (.A1(_04032_),
    .A2(_04096_),
    .B(_03644_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09749_ (.A1(_02298_),
    .A2(_03614_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09750_ (.I(_04077_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09751_ (.I(_03784_),
    .Z(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09752_ (.I(_02254_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09753_ (.I(_04101_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09754_ (.I(_03783_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09755_ (.I(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09756_ (.A1(\as2650.stack[2][2] ),
    .A2(_04102_),
    .B1(_04104_),
    .B2(\as2650.stack[3][2] ),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09757_ (.I(_02470_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09758_ (.I(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09759_ (.I(_02586_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09760_ (.I(_04108_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09761_ (.A1(\as2650.stack[1][2] ),
    .A2(_04107_),
    .B1(_04109_),
    .B2(\as2650.stack[0][2] ),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09762_ (.A1(_04100_),
    .A2(_04105_),
    .A3(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09763_ (.I(_03800_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09764_ (.A1(\as2650.stack[5][2] ),
    .A2(_04107_),
    .B1(_04109_),
    .B2(\as2650.stack[4][2] ),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09765_ (.A1(\as2650.stack[6][2] ),
    .A2(_04102_),
    .B1(_04104_),
    .B2(\as2650.stack[7][2] ),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09766_ (.A1(_04112_),
    .A2(_04113_),
    .A3(_04114_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09767_ (.A1(_03780_),
    .A2(_04111_),
    .A3(_04115_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09768_ (.A1(\as2650.stack[10][2] ),
    .A2(_03998_),
    .B1(_03999_),
    .B2(\as2650.stack[11][2] ),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09769_ (.A1(\as2650.stack[9][2] ),
    .A2(_03995_),
    .B1(_03996_),
    .B2(\as2650.stack[8][2] ),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09770_ (.A1(_04100_),
    .A2(_04117_),
    .A3(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09771_ (.A1(\as2650.stack[13][2] ),
    .A2(_04107_),
    .B1(_04109_),
    .B2(\as2650.stack[12][2] ),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09772_ (.A1(\as2650.stack[14][2] ),
    .A2(_04102_),
    .B1(_04104_),
    .B2(\as2650.stack[15][2] ),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09773_ (.A1(_03801_),
    .A2(_04120_),
    .A3(_04121_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09774_ (.A1(_03812_),
    .A2(_04119_),
    .A3(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09775_ (.A1(_04116_),
    .A2(_04123_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09776_ (.A1(_03434_),
    .A2(_04050_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09777_ (.A1(_04099_),
    .A2(_04124_),
    .B(_04125_),
    .C(_04039_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09778_ (.I(_03686_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09779_ (.A1(_02298_),
    .A2(_04043_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09780_ (.A1(_03687_),
    .A2(_04128_),
    .B(_04079_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09781_ (.A1(_02300_),
    .A2(_04127_),
    .B(_04129_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09782_ (.I(_03709_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09783_ (.A1(_04126_),
    .A2(_04130_),
    .B(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09784_ (.A1(_04098_),
    .A2(_04132_),
    .B(_01688_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09785_ (.A1(_03426_),
    .A2(_03824_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09786_ (.A1(_03969_),
    .A2(_04098_),
    .A3(_04132_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09787_ (.A1(_04096_),
    .A2(_04135_),
    .B(_04087_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09788_ (.A1(_04022_),
    .A2(_04134_),
    .A3(_04136_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09789_ (.A1(_04036_),
    .A2(_04133_),
    .A3(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09790_ (.A1(_03897_),
    .A2(_04095_),
    .B1(_04097_),
    .B2(_04138_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09791_ (.A1(_04030_),
    .A2(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09792_ (.A1(_03081_),
    .A2(_04093_),
    .B(_04140_),
    .C(_04029_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09793_ (.I(_03704_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09794_ (.I(_03666_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09795_ (.I(_04087_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09796_ (.I(_03636_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09797_ (.A1(_02297_),
    .A2(\as2650.PC[3] ),
    .A3(_04043_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09798_ (.A1(_02298_),
    .A2(_04043_),
    .B(\as2650.PC[3] ),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09799_ (.A1(_02309_),
    .A2(_04041_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09800_ (.A1(_04041_),
    .A2(_04145_),
    .A3(_04146_),
    .B(_04147_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09801_ (.I(_03636_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09802_ (.I(_04049_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09803_ (.I(_04150_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09804_ (.A1(_02309_),
    .A2(_04151_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09805_ (.I(_03790_),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09806_ (.A1(\as2650.stack[2][3] ),
    .A2(_04063_),
    .B1(_04153_),
    .B2(\as2650.stack[3][3] ),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09807_ (.A1(\as2650.stack[1][3] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(\as2650.stack[0][3] ),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09808_ (.A1(_04052_),
    .A2(_04154_),
    .A3(_04155_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09809_ (.I(_02472_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09810_ (.I(_02588_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09811_ (.A1(\as2650.stack[5][3] ),
    .A2(_04157_),
    .B1(_04158_),
    .B2(\as2650.stack[4][3] ),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09812_ (.I(_02256_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09813_ (.A1(\as2650.stack[6][3] ),
    .A2(_04160_),
    .B1(_04054_),
    .B2(\as2650.stack[7][3] ),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09814_ (.A1(_04071_),
    .A2(_04159_),
    .A3(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09815_ (.A1(_04051_),
    .A2(_04156_),
    .A3(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09816_ (.I(_03785_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09817_ (.A1(\as2650.stack[10][3] ),
    .A2(_04160_),
    .B1(_04153_),
    .B2(\as2650.stack[11][3] ),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09818_ (.A1(\as2650.stack[9][3] ),
    .A2(_04157_),
    .B1(_04158_),
    .B2(\as2650.stack[8][3] ),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09819_ (.A1(_04164_),
    .A2(_04165_),
    .A3(_04166_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09820_ (.A1(\as2650.stack[13][3] ),
    .A2(_04157_),
    .B1(_04158_),
    .B2(\as2650.stack[12][3] ),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09821_ (.A1(\as2650.stack[14][3] ),
    .A2(_04160_),
    .B1(_04153_),
    .B2(\as2650.stack[15][3] ),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09822_ (.A1(_04071_),
    .A2(_04168_),
    .A3(_04169_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09823_ (.A1(_04003_),
    .A2(_04167_),
    .A3(_04170_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09824_ (.A1(_04163_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09825_ (.A1(_03981_),
    .A2(_04172_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09826_ (.A1(_04149_),
    .A2(_04152_),
    .A3(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09827_ (.A1(_04144_),
    .A2(_04148_),
    .B(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09828_ (.A1(_03738_),
    .A2(_04175_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09829_ (.A1(\as2650.PC[3] ),
    .A2(_03615_),
    .B(_04176_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09830_ (.A1(_04085_),
    .A2(_02309_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09831_ (.A1(_03970_),
    .A2(_04177_),
    .B(_04178_),
    .C(_04143_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09832_ (.A1(_03443_),
    .A2(_04143_),
    .B(_04179_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09833_ (.A1(_04142_),
    .A2(_04180_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09834_ (.A1(_04021_),
    .A2(_03971_),
    .B(_03385_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09835_ (.I(_04182_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09836_ (.A1(_01689_),
    .A2(_04177_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09837_ (.A1(_04181_),
    .A2(_04183_),
    .A3(_04184_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09838_ (.I(_04178_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09839_ (.A1(_03708_),
    .A2(_03971_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09840_ (.A1(_03843_),
    .A2(_03845_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09841_ (.A1(_03770_),
    .A2(_04188_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09842_ (.A1(_03843_),
    .A2(_03845_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09843_ (.A1(_04186_),
    .A2(_04187_),
    .B1(_04189_),
    .B2(_04190_),
    .C(_03867_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09844_ (.A1(_03749_),
    .A2(_04141_),
    .B1(_04185_),
    .B2(_04191_),
    .C(_03520_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09845_ (.A1(_03970_),
    .A2(_02326_),
    .B(_04032_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09846_ (.A1(_02321_),
    .A2(_04145_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09847_ (.A1(_02325_),
    .A2(_04040_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09848_ (.A1(_04046_),
    .A2(_04193_),
    .B(_04194_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09849_ (.I(_02255_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09850_ (.I(_03789_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09851_ (.A1(\as2650.stack[2][4] ),
    .A2(_04196_),
    .B1(_04197_),
    .B2(\as2650.stack[3][4] ),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09852_ (.I(_02471_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09853_ (.I(_02587_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09854_ (.A1(\as2650.stack[1][4] ),
    .A2(_04199_),
    .B1(_04200_),
    .B2(\as2650.stack[0][4] ),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09855_ (.A1(_03785_),
    .A2(_04198_),
    .A3(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09856_ (.I(_02471_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09857_ (.I(_02587_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09858_ (.A1(\as2650.stack[5][4] ),
    .A2(_04203_),
    .B1(_04204_),
    .B2(\as2650.stack[4][4] ),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09859_ (.I(_02255_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09860_ (.I(_03789_),
    .Z(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09861_ (.A1(\as2650.stack[6][4] ),
    .A2(_04206_),
    .B1(_04207_),
    .B2(\as2650.stack[7][4] ),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09862_ (.A1(_04007_),
    .A2(_04205_),
    .A3(_04208_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09863_ (.A1(_03779_),
    .A2(_04202_),
    .A3(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09864_ (.A1(\as2650.stack[10][4] ),
    .A2(_04196_),
    .B1(_04197_),
    .B2(\as2650.stack[11][4] ),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09865_ (.A1(\as2650.stack[9][4] ),
    .A2(_04199_),
    .B1(_04200_),
    .B2(\as2650.stack[8][4] ),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09866_ (.A1(_04100_),
    .A2(_04211_),
    .A3(_04212_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09867_ (.A1(\as2650.stack[13][4] ),
    .A2(_04203_),
    .B1(_04204_),
    .B2(\as2650.stack[12][4] ),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09868_ (.A1(\as2650.stack[14][4] ),
    .A2(_04206_),
    .B1(_04207_),
    .B2(\as2650.stack[15][4] ),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09869_ (.A1(_04112_),
    .A2(_04214_),
    .A3(_04215_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09870_ (.A1(_03812_),
    .A2(_04213_),
    .A3(_04216_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09871_ (.A1(_04210_),
    .A2(_04217_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09872_ (.A1(_02325_),
    .A2(_04150_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09873_ (.A1(_04077_),
    .A2(_04218_),
    .B(_04219_),
    .C(_04038_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09874_ (.A1(_04079_),
    .A2(_04195_),
    .B(_04220_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09875_ (.A1(_03772_),
    .A2(_04221_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09876_ (.A1(_02321_),
    .A2(_03614_),
    .B(_04222_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09877_ (.A1(_01688_),
    .A2(_04223_),
    .B(_03973_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09878_ (.A1(_03969_),
    .A2(_04223_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09879_ (.A1(_04021_),
    .A2(_02326_),
    .B(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09880_ (.I(_03823_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09881_ (.A1(_03172_),
    .A2(_03406_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09882_ (.A1(_03441_),
    .A2(_03465_),
    .B(_04227_),
    .C(_04228_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09883_ (.A1(_03975_),
    .A2(_04226_),
    .B(_04229_),
    .C(_04022_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09884_ (.A1(_04224_),
    .A2(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09885_ (.A1(_03968_),
    .A2(_04192_),
    .B(_04231_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09886_ (.A1(net200),
    .A2(_03854_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09887_ (.A1(_03469_),
    .A2(_04233_),
    .A3(_03847_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09888_ (.A1(_03925_),
    .A2(_04234_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09889_ (.A1(_04232_),
    .A2(_04235_),
    .B(_03765_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09890_ (.A1(_03753_),
    .A2(_04093_),
    .B(_04236_),
    .C(_04029_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09891_ (.I(_03737_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09892_ (.I(_04038_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09893_ (.I(_04040_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _09894_ (.A1(_02320_),
    .A2(_02337_),
    .A3(_04145_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09895_ (.A1(_02321_),
    .A2(_04145_),
    .B(_02337_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09896_ (.A1(_02341_),
    .A2(_04046_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _09897_ (.A1(_04239_),
    .A2(_04240_),
    .A3(_04241_),
    .B(_04242_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09898_ (.A1(_02342_),
    .A2(_04150_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09899_ (.A1(\as2650.stack[2][5] ),
    .A2(_04206_),
    .B1(_04207_),
    .B2(\as2650.stack[3][5] ),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09900_ (.A1(\as2650.stack[1][5] ),
    .A2(_04203_),
    .B1(_04204_),
    .B2(\as2650.stack[0][5] ),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09901_ (.A1(_03785_),
    .A2(_04245_),
    .A3(_04246_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09902_ (.A1(\as2650.stack[5][5] ),
    .A2(_04203_),
    .B1(_04204_),
    .B2(\as2650.stack[4][5] ),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09903_ (.A1(\as2650.stack[6][5] ),
    .A2(_04206_),
    .B1(_04207_),
    .B2(\as2650.stack[7][5] ),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09904_ (.A1(_04112_),
    .A2(_04248_),
    .A3(_04249_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09905_ (.A1(_03779_),
    .A2(_04247_),
    .A3(_04250_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09906_ (.A1(\as2650.stack[10][5] ),
    .A2(_04196_),
    .B1(_04197_),
    .B2(\as2650.stack[11][5] ),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09907_ (.A1(\as2650.stack[9][5] ),
    .A2(_04199_),
    .B1(_04200_),
    .B2(\as2650.stack[8][5] ),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09908_ (.A1(_04100_),
    .A2(_04252_),
    .A3(_04253_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09909_ (.A1(\as2650.stack[13][5] ),
    .A2(_04199_),
    .B1(_04200_),
    .B2(\as2650.stack[12][5] ),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09910_ (.A1(\as2650.stack[14][5] ),
    .A2(_04196_),
    .B1(_04197_),
    .B2(\as2650.stack[15][5] ),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09911_ (.A1(_04112_),
    .A2(_04255_),
    .A3(_04256_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09912_ (.A1(_03812_),
    .A2(_04254_),
    .A3(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09913_ (.A1(_04251_),
    .A2(_04258_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09914_ (.A1(_03773_),
    .A2(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09915_ (.A1(_04079_),
    .A2(_04244_),
    .A3(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09916_ (.A1(_04238_),
    .A2(_04243_),
    .B(_04261_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09917_ (.A1(_03772_),
    .A2(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09918_ (.A1(_02337_),
    .A2(_04237_),
    .B(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09919_ (.A1(_03969_),
    .A2(_02342_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09920_ (.A1(_04085_),
    .A2(_04264_),
    .B(_04265_),
    .C(_04087_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09921_ (.A1(_03480_),
    .A2(_03875_),
    .B(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09922_ (.A1(_03903_),
    .A2(_04267_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09923_ (.A1(_04037_),
    .A2(_04264_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09924_ (.A1(_04182_),
    .A2(_04268_),
    .A3(_04269_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09925_ (.A1(_03849_),
    .A2(_03852_),
    .B(_03770_),
    .ZN(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09926_ (.A1(_03849_),
    .A2(_03852_),
    .B(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09927_ (.A1(_03970_),
    .A2(_02342_),
    .A3(_04187_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09928_ (.A1(_03733_),
    .A2(_04270_),
    .A3(_04272_),
    .A4(_04273_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09929_ (.I(_03963_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09930_ (.A1(_03756_),
    .A2(_04093_),
    .B(_04274_),
    .C(_04275_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09931_ (.I(_03561_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09932_ (.A1(\as2650.stack[2][6] ),
    .A2(_04101_),
    .B1(_04103_),
    .B2(\as2650.stack[3][6] ),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09933_ (.A1(\as2650.stack[1][6] ),
    .A2(_04106_),
    .B1(_04108_),
    .B2(\as2650.stack[0][6] ),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09934_ (.A1(_03982_),
    .A2(_04277_),
    .A3(_04278_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09935_ (.A1(\as2650.stack[5][6] ),
    .A2(_04106_),
    .B1(_04108_),
    .B2(\as2650.stack[4][6] ),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09936_ (.A1(\as2650.stack[6][6] ),
    .A2(_04101_),
    .B1(_04103_),
    .B2(\as2650.stack[7][6] ),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09937_ (.A1(_03800_),
    .A2(_04280_),
    .A3(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09938_ (.A1(_03778_),
    .A2(_04279_),
    .A3(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09939_ (.A1(\as2650.stack[10][6] ),
    .A2(_03984_),
    .B1(_03986_),
    .B2(\as2650.stack[11][6] ),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09940_ (.A1(\as2650.stack[9][6] ),
    .A2(_03989_),
    .B1(_04108_),
    .B2(\as2650.stack[8][6] ),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09941_ (.A1(_03982_),
    .A2(_04284_),
    .A3(_04285_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09942_ (.A1(\as2650.stack[13][6] ),
    .A2(_04106_),
    .B1(_03991_),
    .B2(\as2650.stack[12][6] ),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09943_ (.A1(\as2650.stack[14][6] ),
    .A2(_04101_),
    .B1(_04103_),
    .B2(\as2650.stack[15][6] ),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09944_ (.A1(_03800_),
    .A2(_04287_),
    .A3(_04288_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09945_ (.A1(_03811_),
    .A2(_04286_),
    .A3(_04289_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09946_ (.A1(_04283_),
    .A2(_04290_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09947_ (.I(_04291_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09948_ (.A1(_03981_),
    .A2(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09949_ (.A1(_02357_),
    .A2(_03774_),
    .B(_04293_),
    .C(_04144_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09950_ (.A1(_02353_),
    .A2(_04240_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09951_ (.A1(_04127_),
    .A2(_04295_),
    .B(_04039_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09952_ (.A1(_02357_),
    .A2(_03688_),
    .B(_04296_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09953_ (.A1(_03738_),
    .A2(_04294_),
    .A3(_04297_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09954_ (.A1(_02353_),
    .A2(_03615_),
    .B(_04298_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09955_ (.A1(_04085_),
    .A2(_02357_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09956_ (.A1(_04021_),
    .A2(_04299_),
    .B(_04300_),
    .C(_03875_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09957_ (.I(_04227_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09958_ (.A1(_03440_),
    .A2(_03496_),
    .B(_03487_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09959_ (.A1(_04302_),
    .A2(_04303_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09960_ (.A1(_04301_),
    .A2(_04304_),
    .B(_04037_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09961_ (.A1(_04276_),
    .A2(_04299_),
    .B(_04305_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09962_ (.A1(_04183_),
    .A2(_04306_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09963_ (.I(_04300_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09964_ (.A1(net203),
    .A2(_03854_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09965_ (.A1(_03500_),
    .A2(_04309_),
    .A3(_03853_),
    .Z(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09966_ (.A1(_04187_),
    .A2(_04308_),
    .B1(_04310_),
    .B2(_03870_),
    .C(_03867_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _09967_ (.A1(_03758_),
    .A2(_04141_),
    .B1(_04307_),
    .B2(_04311_),
    .C(_03520_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09968_ (.A1(_03440_),
    .A2(_03511_),
    .B(_03488_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09969_ (.I(_04050_),
    .Z(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09970_ (.I(_03983_),
    .Z(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09971_ (.I(_03998_),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09972_ (.I(_03999_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09973_ (.A1(\as2650.stack[2][7] ),
    .A2(_04315_),
    .B1(_04316_),
    .B2(\as2650.stack[3][7] ),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09974_ (.I(_03995_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09975_ (.I(_03996_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09976_ (.A1(\as2650.stack[1][7] ),
    .A2(_04318_),
    .B1(_04319_),
    .B2(\as2650.stack[0][7] ),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09977_ (.A1(_04314_),
    .A2(_04317_),
    .A3(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09978_ (.I(_03801_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09979_ (.A1(\as2650.stack[5][7] ),
    .A2(_04318_),
    .B1(_04319_),
    .B2(\as2650.stack[4][7] ),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09980_ (.A1(\as2650.stack[6][7] ),
    .A2(_04315_),
    .B1(_04316_),
    .B2(\as2650.stack[7][7] ),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09981_ (.A1(_04322_),
    .A2(_04323_),
    .A3(_04324_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09982_ (.A1(_03781_),
    .A2(_04321_),
    .A3(_04325_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09983_ (.I(_03998_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09984_ (.I(_03999_),
    .Z(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09985_ (.A1(\as2650.stack[10][7] ),
    .A2(_04327_),
    .B1(_04328_),
    .B2(\as2650.stack[11][7] ),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09986_ (.I(_03995_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09987_ (.I(_03996_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09988_ (.A1(\as2650.stack[9][7] ),
    .A2(_04330_),
    .B1(_04331_),
    .B2(\as2650.stack[8][7] ),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09989_ (.A1(_04314_),
    .A2(_04329_),
    .A3(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09990_ (.A1(\as2650.stack[13][7] ),
    .A2(_04318_),
    .B1(_04319_),
    .B2(\as2650.stack[12][7] ),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09991_ (.A1(\as2650.stack[14][7] ),
    .A2(_04315_),
    .B1(_04316_),
    .B2(\as2650.stack[15][7] ),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09992_ (.A1(_04322_),
    .A2(_04334_),
    .A3(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09993_ (.A1(_03813_),
    .A2(_04333_),
    .A3(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _09994_ (.A1(_04326_),
    .A2(_04337_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09995_ (.A1(_03524_),
    .A2(_04099_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09996_ (.A1(_04313_),
    .A2(_04338_),
    .B(_04339_),
    .C(_03637_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09997_ (.A1(_02353_),
    .A2(_04240_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09998_ (.A1(_02381_),
    .A2(_04341_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09999_ (.A1(_04127_),
    .A2(_04342_),
    .B(_04144_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10000_ (.A1(_02369_),
    .A2(_03688_),
    .B(_04343_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10001_ (.A1(_04340_),
    .A2(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10002_ (.A1(_02367_),
    .A2(_04017_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10003_ (.A1(_04017_),
    .A2(_04345_),
    .B(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10004_ (.I(_00953_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10005_ (.A1(_04348_),
    .A2(_02369_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10006_ (.A1(_03974_),
    .A2(_04347_),
    .B(_04349_),
    .C(_04302_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10007_ (.A1(_04302_),
    .A2(_04312_),
    .B(_04350_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10008_ (.I(_04017_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10009_ (.A1(_04352_),
    .A2(_04345_),
    .B(_04346_),
    .C(_04276_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10010_ (.A1(_01689_),
    .A2(_04351_),
    .B(_04353_),
    .C(_04183_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10011_ (.A1(_03856_),
    .A2(_03859_),
    .B(_03869_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10012_ (.A1(_03856_),
    .A2(_03859_),
    .B(_04355_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10013_ (.A1(_04187_),
    .A2(_04349_),
    .B(_04356_),
    .C(_03704_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10014_ (.A1(_03762_),
    .A2(_04141_),
    .B1(_04354_),
    .B2(_04357_),
    .C(_03520_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10015_ (.A1(_03828_),
    .A2(_03861_),
    .Z(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10016_ (.I(_03971_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10017_ (.A1(_04020_),
    .A2(_02384_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10018_ (.A1(_04359_),
    .A2(_04360_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10019_ (.A1(_03440_),
    .A2(_03528_),
    .B(_03487_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10020_ (.A1(_02352_),
    .A2(_02367_),
    .A3(_04240_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10021_ (.A1(_02385_),
    .A2(_04363_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10022_ (.A1(_02385_),
    .A2(_04363_),
    .B(_03686_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10023_ (.A1(_02384_),
    .A2(_04239_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10024_ (.A1(_04364_),
    .A2(_04365_),
    .B(_04366_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10025_ (.I(_02256_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10026_ (.I(_03790_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10027_ (.A1(\as2650.stack[2][8] ),
    .A2(_04368_),
    .B1(_04369_),
    .B2(\as2650.stack[3][8] ),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10028_ (.I(_02472_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10029_ (.I(_02588_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10030_ (.A1(\as2650.stack[1][8] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\as2650.stack[0][8] ),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10031_ (.A1(_04164_),
    .A2(_04370_),
    .A3(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10032_ (.I(_04007_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10033_ (.A1(\as2650.stack[5][8] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\as2650.stack[4][8] ),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10034_ (.A1(\as2650.stack[6][8] ),
    .A2(_04368_),
    .B1(_04369_),
    .B2(\as2650.stack[7][8] ),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10035_ (.A1(_04375_),
    .A2(_04376_),
    .A3(_04377_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10036_ (.A1(_04051_),
    .A2(_04374_),
    .A3(_04378_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10037_ (.I(_03811_),
    .Z(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10038_ (.A1(\as2650.stack[10][8] ),
    .A2(_04368_),
    .B1(_04369_),
    .B2(\as2650.stack[11][8] ),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10039_ (.A1(\as2650.stack[9][8] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\as2650.stack[8][8] ),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10040_ (.A1(_03786_),
    .A2(_04381_),
    .A3(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10041_ (.A1(\as2650.stack[13][8] ),
    .A2(_04371_),
    .B1(_04372_),
    .B2(\as2650.stack[12][8] ),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10042_ (.A1(\as2650.stack[14][8] ),
    .A2(_04368_),
    .B1(_04369_),
    .B2(\as2650.stack[15][8] ),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10043_ (.A1(_04375_),
    .A2(_04384_),
    .A3(_04385_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10044_ (.A1(_04380_),
    .A2(_04383_),
    .A3(_04386_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10045_ (.A1(_04379_),
    .A2(_04387_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10046_ (.A1(_02384_),
    .A2(_04050_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10047_ (.A1(_04151_),
    .A2(_04388_),
    .B(_04389_),
    .C(_04238_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10048_ (.A1(_04144_),
    .A2(_04367_),
    .B(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10049_ (.A1(_02380_),
    .A2(_04131_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10050_ (.A1(_03710_),
    .A2(_04391_),
    .B(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10051_ (.A1(_04348_),
    .A2(_04393_),
    .B(_04360_),
    .C(_04227_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10052_ (.A1(_04302_),
    .A2(_04362_),
    .B(_04394_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10053_ (.A1(_03711_),
    .A2(_04391_),
    .B(_04392_),
    .C(_01688_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10054_ (.I(_04036_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10055_ (.A1(_04276_),
    .A2(_04395_),
    .B(_04396_),
    .C(_04397_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10056_ (.A1(_03968_),
    .A2(_04361_),
    .B(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10057_ (.A1(_03771_),
    .A2(_04358_),
    .B(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10058_ (.I(_01448_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10059_ (.A1(\as2650.instruction_args_latch[8] ),
    .A2(_03733_),
    .B(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10060_ (.A1(_03929_),
    .A2(_04400_),
    .B(_04402_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10061_ (.A1(_03828_),
    .A2(_03861_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10062_ (.A1(_03404_),
    .A2(_04403_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10063_ (.A1(_03925_),
    .A2(_04404_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10064_ (.A1(_04020_),
    .A2(_02399_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10065_ (.A1(_04032_),
    .A2(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10066_ (.A1(_02380_),
    .A2(_02396_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10067_ (.A1(_04363_),
    .A2(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10068_ (.A1(_02399_),
    .A2(_04046_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10069_ (.A1(_04239_),
    .A2(_04409_),
    .B(_04410_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10070_ (.A1(\as2650.stack[2][9] ),
    .A2(_04053_),
    .B1(_04064_),
    .B2(\as2650.stack[3][9] ),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10071_ (.A1(\as2650.stack[1][9] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[0][9] ),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10072_ (.A1(_03983_),
    .A2(_04412_),
    .A3(_04413_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10073_ (.A1(\as2650.stack[5][9] ),
    .A2(_03990_),
    .B1(_03992_),
    .B2(\as2650.stack[4][9] ),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10074_ (.A1(\as2650.stack[6][9] ),
    .A2(_03985_),
    .B1(_03987_),
    .B2(\as2650.stack[7][9] ),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10075_ (.A1(_04008_),
    .A2(_04415_),
    .A3(_04416_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10076_ (.A1(_03780_),
    .A2(_04414_),
    .A3(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10077_ (.A1(\as2650.stack[10][9] ),
    .A2(_04053_),
    .B1(_04064_),
    .B2(\as2650.stack[11][9] ),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10078_ (.A1(\as2650.stack[9][9] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[8][9] ),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10079_ (.A1(_04052_),
    .A2(_04419_),
    .A3(_04420_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10080_ (.A1(\as2650.stack[13][9] ),
    .A2(_04056_),
    .B1(_04057_),
    .B2(\as2650.stack[12][9] ),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10081_ (.A1(\as2650.stack[14][9] ),
    .A2(_04053_),
    .B1(_04064_),
    .B2(\as2650.stack[15][9] ),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10082_ (.A1(_04008_),
    .A2(_04422_),
    .A3(_04423_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10083_ (.A1(_04003_),
    .A2(_04421_),
    .A3(_04424_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10084_ (.A1(_04418_),
    .A2(_04425_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10085_ (.A1(_02398_),
    .A2(_04150_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10086_ (.A1(_04077_),
    .A2(_04426_),
    .B(_04427_),
    .C(_03636_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10087_ (.A1(_04039_),
    .A2(_04411_),
    .B(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10088_ (.A1(_03737_),
    .A2(_04365_),
    .B(_02396_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10089_ (.A1(_03772_),
    .A2(_04429_),
    .B(_04430_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10090_ (.A1(_03369_),
    .A2(_04227_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10091_ (.A1(_04033_),
    .A2(_04431_),
    .B(_04406_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10092_ (.A1(_03541_),
    .A2(_04432_),
    .B1(_04433_),
    .B2(_03824_),
    .C(_03666_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10093_ (.A1(_03903_),
    .A2(_04431_),
    .B(_04434_),
    .C(_04036_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10094_ (.A1(_03968_),
    .A2(_04407_),
    .B(_04435_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10095_ (.A1(_04405_),
    .A2(_04436_),
    .B(_03704_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10096_ (.A1(_01151_),
    .A2(_04093_),
    .B(_04437_),
    .C(_04275_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10097_ (.I(_04022_),
    .Z(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10098_ (.A1(\as2650.stack[2][10] ),
    .A2(_04315_),
    .B1(_04316_),
    .B2(\as2650.stack[3][10] ),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10099_ (.A1(\as2650.stack[1][10] ),
    .A2(_04318_),
    .B1(_04319_),
    .B2(\as2650.stack[0][10] ),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10100_ (.A1(_04314_),
    .A2(_04439_),
    .A3(_04440_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10101_ (.A1(\as2650.stack[5][10] ),
    .A2(_04330_),
    .B1(_04331_),
    .B2(\as2650.stack[4][10] ),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10102_ (.A1(\as2650.stack[6][10] ),
    .A2(_04327_),
    .B1(_04328_),
    .B2(\as2650.stack[7][10] ),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10103_ (.A1(_04322_),
    .A2(_04442_),
    .A3(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10104_ (.A1(_03781_),
    .A2(_04441_),
    .A3(_04444_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10105_ (.A1(\as2650.stack[10][10] ),
    .A2(_04327_),
    .B1(_04328_),
    .B2(\as2650.stack[11][10] ),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10106_ (.A1(\as2650.stack[9][10] ),
    .A2(_04330_),
    .B1(_04331_),
    .B2(\as2650.stack[8][10] ),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10107_ (.A1(_04314_),
    .A2(_04446_),
    .A3(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10108_ (.A1(\as2650.stack[13][10] ),
    .A2(_04330_),
    .B1(_04331_),
    .B2(\as2650.stack[12][10] ),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10109_ (.A1(\as2650.stack[14][10] ),
    .A2(_04327_),
    .B1(_04328_),
    .B2(\as2650.stack[15][10] ),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10110_ (.A1(_03802_),
    .A2(_04449_),
    .A3(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10111_ (.A1(_04380_),
    .A2(_04448_),
    .A3(_04451_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10112_ (.A1(_03981_),
    .A2(_04445_),
    .A3(_04452_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10113_ (.A1(_02414_),
    .A2(_03774_),
    .B(_04453_),
    .C(_04149_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10114_ (.A1(_02410_),
    .A2(_04409_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10115_ (.A1(_03687_),
    .A2(_04455_),
    .B(_04238_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10116_ (.A1(_02414_),
    .A2(_04127_),
    .B(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10117_ (.A1(_04237_),
    .A2(_04454_),
    .A3(_04457_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10118_ (.A1(_02409_),
    .A2(_03738_),
    .B(_04458_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10119_ (.A1(_04033_),
    .A2(_02414_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10120_ (.A1(_03974_),
    .A2(_04459_),
    .B(_04460_),
    .C(_03975_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10121_ (.A1(_03555_),
    .A2(_04432_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10122_ (.A1(_04461_),
    .A2(_04462_),
    .B(_03903_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10123_ (.A1(_04438_),
    .A2(_04459_),
    .B(_04463_),
    .C(_04397_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10124_ (.A1(_04359_),
    .A2(_04460_),
    .B(_03642_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10125_ (.A1(_03403_),
    .A2(_04403_),
    .B(_03420_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10126_ (.A1(_03862_),
    .A2(_03771_),
    .A3(_04466_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10127_ (.A1(_04464_),
    .A2(_04465_),
    .B(_04467_),
    .C(_03927_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10128_ (.A1(_03418_),
    .A2(_03929_),
    .B(_03930_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10129_ (.A1(_04468_),
    .A2(_04469_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10130_ (.I(\as2650.instruction_args_latch[11] ),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10131_ (.A1(_02409_),
    .A2(_04409_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10132_ (.A1(_03688_),
    .A2(_04471_),
    .B(_04131_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10133_ (.A1(\as2650.stack[2][11] ),
    .A2(_02257_),
    .B1(_03791_),
    .B2(\as2650.stack[3][11] ),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10134_ (.A1(\as2650.stack[1][11] ),
    .A2(_02473_),
    .B1(_02589_),
    .B2(\as2650.stack[0][11] ),
    .ZN(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10135_ (.A1(_04164_),
    .A2(_04473_),
    .A3(_04474_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10136_ (.A1(\as2650.stack[5][11] ),
    .A2(_04157_),
    .B1(_04158_),
    .B2(\as2650.stack[4][11] ),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10137_ (.A1(\as2650.stack[6][11] ),
    .A2(_04160_),
    .B1(_04153_),
    .B2(\as2650.stack[7][11] ),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10138_ (.A1(_04071_),
    .A2(_04476_),
    .A3(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10139_ (.A1(_04051_),
    .A2(_04475_),
    .A3(_04478_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10140_ (.A1(\as2650.stack[10][11] ),
    .A2(_02257_),
    .B1(_03791_),
    .B2(\as2650.stack[11][11] ),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10141_ (.A1(\as2650.stack[9][11] ),
    .A2(_02473_),
    .B1(_02589_),
    .B2(\as2650.stack[8][11] ),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10142_ (.A1(_04164_),
    .A2(_04480_),
    .A3(_04481_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10143_ (.A1(\as2650.stack[13][11] ),
    .A2(_02473_),
    .B1(_02589_),
    .B2(\as2650.stack[12][11] ),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10144_ (.A1(\as2650.stack[14][11] ),
    .A2(_02257_),
    .B1(_03791_),
    .B2(\as2650.stack[15][11] ),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10145_ (.A1(_04375_),
    .A2(_04483_),
    .A3(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10146_ (.A1(_04380_),
    .A2(_04482_),
    .A3(_04485_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10147_ (.A1(_04479_),
    .A2(_04486_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10148_ (.A1(_04151_),
    .A2(_04487_),
    .B(_04238_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10149_ (.A1(_02427_),
    .A2(_04099_),
    .B(_04488_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10150_ (.A1(_02409_),
    .A2(_02424_),
    .A3(_04409_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10151_ (.A1(_03686_),
    .A2(_04490_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10152_ (.A1(_02427_),
    .A2(_04041_),
    .B(_04149_),
    .C(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10153_ (.A1(_04489_),
    .A2(_04492_),
    .B(_04237_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10154_ (.A1(_02424_),
    .A2(_04472_),
    .B(_04493_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10155_ (.A1(_04348_),
    .A2(_02427_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10156_ (.A1(_03974_),
    .A2(_04494_),
    .B(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10157_ (.A1(_03569_),
    .A2(_03876_),
    .B1(_04496_),
    .B2(_04143_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10158_ (.A1(_04276_),
    .A2(_04497_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10159_ (.A1(_04438_),
    .A2(_04494_),
    .B(_04397_),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10160_ (.A1(_04359_),
    .A2(_04495_),
    .B(_03642_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10161_ (.A1(_04498_),
    .A2(_04499_),
    .B(_04500_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10162_ (.A1(_03560_),
    .A2(_03862_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10163_ (.A1(_03560_),
    .A2(_03862_),
    .B(_03897_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10164_ (.I(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10165_ (.A1(_04502_),
    .A2(_04504_),
    .B(_04030_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10166_ (.A1(_04470_),
    .A2(_04141_),
    .B1(_04501_),
    .B2(_04505_),
    .C(_01460_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10167_ (.I(_04102_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10168_ (.I(_04104_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10169_ (.A1(\as2650.stack[2][12] ),
    .A2(_04506_),
    .B1(_04507_),
    .B2(\as2650.stack[3][12] ),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10170_ (.I(_04107_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10171_ (.I(_04109_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10172_ (.A1(\as2650.stack[1][12] ),
    .A2(_04509_),
    .B1(_04510_),
    .B2(\as2650.stack[0][12] ),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10173_ (.A1(_03786_),
    .A2(_04508_),
    .A3(_04511_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10174_ (.A1(\as2650.stack[5][12] ),
    .A2(_04509_),
    .B1(_04510_),
    .B2(\as2650.stack[4][12] ),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10175_ (.A1(\as2650.stack[6][12] ),
    .A2(_04506_),
    .B1(_04507_),
    .B2(\as2650.stack[7][12] ),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10176_ (.A1(_04375_),
    .A2(_04513_),
    .A3(_04514_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10177_ (.A1(_03781_),
    .A2(_04512_),
    .A3(_04515_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10178_ (.A1(\as2650.stack[10][12] ),
    .A2(_04506_),
    .B1(_04507_),
    .B2(\as2650.stack[11][12] ),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10179_ (.A1(\as2650.stack[9][12] ),
    .A2(_04509_),
    .B1(_04510_),
    .B2(\as2650.stack[8][12] ),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10180_ (.A1(_03786_),
    .A2(_04517_),
    .A3(_04518_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10181_ (.A1(\as2650.stack[13][12] ),
    .A2(_04509_),
    .B1(_04510_),
    .B2(\as2650.stack[12][12] ),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10182_ (.A1(\as2650.stack[14][12] ),
    .A2(_04506_),
    .B1(_04507_),
    .B2(\as2650.stack[15][12] ),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10183_ (.A1(_04322_),
    .A2(_04520_),
    .A3(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10184_ (.A1(_04380_),
    .A2(_04519_),
    .A3(_04522_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10185_ (.A1(_04516_),
    .A2(_04523_),
    .Z(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10186_ (.A1(_02438_),
    .A2(_04151_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10187_ (.A1(_04099_),
    .A2(_04524_),
    .B(_04525_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10188_ (.A1(_02437_),
    .A2(_04239_),
    .B(_04491_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10189_ (.A1(_02436_),
    .A2(_04527_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10190_ (.A1(_02436_),
    .A2(_04527_),
    .B(_04149_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10191_ (.A1(_03637_),
    .A2(_04526_),
    .B1(_04528_),
    .B2(_04529_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10192_ (.A1(_02436_),
    .A2(_04131_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10193_ (.A1(_03710_),
    .A2(_04530_),
    .B(_04531_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10194_ (.I0(_02439_),
    .I1(_04532_),
    .S(_04348_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10195_ (.A1(_03575_),
    .A2(_03876_),
    .B1(_04533_),
    .B2(_04143_),
    .C(_04037_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10196_ (.A1(_04438_),
    .A2(_04532_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10197_ (.A1(_04534_),
    .A2(_04535_),
    .B(_04183_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10198_ (.A1(_03461_),
    .A2(_04502_),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10199_ (.A1(_02439_),
    .A2(_04359_),
    .A3(_04397_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10200_ (.A1(_03870_),
    .A2(_04537_),
    .B(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10201_ (.A1(_04536_),
    .A2(_04539_),
    .B(_03927_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10202_ (.A1(\as2650.instruction_args_latch[12] ),
    .A2(_03929_),
    .B(_03930_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10203_ (.A1(_04540_),
    .A2(_04541_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10204_ (.I(_02875_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10205_ (.I(_04542_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10206_ (.I(_04543_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10207_ (.I(_03665_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10208_ (.A1(_02834_),
    .A2(_02955_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10209_ (.I(_04546_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10210_ (.A1(_03630_),
    .A2(_03943_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10211_ (.A1(_01527_),
    .A2(_04548_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10212_ (.A1(_02215_),
    .A2(_01416_),
    .A3(_01393_),
    .A4(_02200_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10213_ (.A1(_02877_),
    .A2(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10214_ (.A1(_02834_),
    .A2(_02874_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10215_ (.I(_04552_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10216_ (.A1(_04549_),
    .A2(_04551_),
    .A3(_04553_),
    .Z(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10217_ (.A1(_03709_),
    .A2(_02878_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10218_ (.A1(_02915_),
    .A2(_00794_),
    .A3(_01524_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10219_ (.A1(_00890_),
    .A2(_01526_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10220_ (.I(_04557_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10221_ (.I(_01421_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10222_ (.A1(_04559_),
    .A2(_01399_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10223_ (.A1(_02229_),
    .A2(_04550_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10224_ (.A1(_02229_),
    .A2(_04558_),
    .B(_04560_),
    .C(_04561_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10225_ (.A1(_02233_),
    .A2(_03632_),
    .A3(_04556_),
    .A4(_04562_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10226_ (.A1(_03689_),
    .A2(_04555_),
    .A3(_04563_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10227_ (.I(_04564_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10228_ (.A1(_03184_),
    .A2(_04547_),
    .B(_04554_),
    .C(_04565_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10229_ (.A1(_02877_),
    .A2(_04557_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10230_ (.I(_04567_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10231_ (.A1(_04554_),
    .A2(_04567_),
    .Z(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10232_ (.A1(_01393_),
    .A2(_02875_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10233_ (.I(_04570_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10234_ (.I(_02915_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10235_ (.A1(_03281_),
    .A2(_03289_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10236_ (.A1(_03280_),
    .A2(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10237_ (.I(_03278_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10238_ (.A1(_04575_),
    .A2(_03279_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10239_ (.A1(_03286_),
    .A2(_04576_),
    .B(_03235_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10240_ (.I(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10241_ (.A1(_02227_),
    .A2(_04572_),
    .B1(_03197_),
    .B2(_04574_),
    .C(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10242_ (.I(_03298_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10243_ (.I(_02937_),
    .Z(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10244_ (.A1(_03251_),
    .A2(_04581_),
    .B(_01811_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10245_ (.A1(_01811_),
    .A2(_02187_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10246_ (.A1(_02883_),
    .A2(_04582_),
    .B1(_04583_),
    .B2(_04581_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10247_ (.A1(_02227_),
    .A2(_04580_),
    .B(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10248_ (.A1(_02197_),
    .A2(_01398_),
    .A3(_02840_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10249_ (.A1(_02820_),
    .A2(_04586_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10250_ (.I(_04587_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10251_ (.I(_04588_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10252_ (.A1(net180),
    .A2(_04588_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10253_ (.A1(_01470_),
    .A2(_04589_),
    .B(_04590_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10254_ (.A1(_04581_),
    .A2(_02883_),
    .A3(_04591_),
    .B(_04571_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10255_ (.A1(_04571_),
    .A2(_04579_),
    .B1(_04585_),
    .B2(_04592_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10256_ (.A1(_04569_),
    .A2(_04593_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10257_ (.A1(_04013_),
    .A2(_04568_),
    .B(_04594_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10258_ (.A1(_02228_),
    .A2(_04566_),
    .B1(_04595_),
    .B2(_04565_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10259_ (.A1(_02215_),
    .A2(_02870_),
    .A3(_02843_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10260_ (.I(_04597_),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10261_ (.I(_04598_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10262_ (.I(_02195_),
    .Z(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10263_ (.I(_04600_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10264_ (.I(_04601_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10265_ (.A1(_04602_),
    .A2(_04598_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10266_ (.I(_03729_),
    .Z(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10267_ (.A1(_04544_),
    .A2(_04599_),
    .B(_04603_),
    .C(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10268_ (.I(_02197_),
    .Z(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10269_ (.I(_04606_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10270_ (.I(_04607_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10271_ (.I(_02895_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10272_ (.A1(_02228_),
    .A2(_04609_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10273_ (.A1(_04608_),
    .A2(_04609_),
    .B(_04610_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10274_ (.I(_02821_),
    .Z(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10275_ (.A1(_04612_),
    .A2(_04597_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10276_ (.A1(_04544_),
    .A2(_04579_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10277_ (.A1(_04611_),
    .A2(_04613_),
    .B(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10278_ (.A1(_04596_),
    .A2(_04605_),
    .B1(_04615_),
    .B2(_04604_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10279_ (.A1(_04544_),
    .A2(_04545_),
    .B(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10280_ (.A1(_02958_),
    .A2(_04614_),
    .B(_03930_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10281_ (.A1(_04617_),
    .A2(_04618_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10282_ (.A1(_02160_),
    .A2(_00730_),
    .A3(_03631_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10283_ (.I(_04619_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10284_ (.I(_03729_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10285_ (.A1(_04612_),
    .A2(_04621_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10286_ (.A1(_04620_),
    .A2(_04622_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10287_ (.I(_04623_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10288_ (.I(_04606_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10289_ (.A1(_02972_),
    .A2(_04625_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10290_ (.A1(_02272_),
    .A2(_03744_),
    .B(_04626_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10291_ (.I(_04237_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10292_ (.I(_04628_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10293_ (.A1(_00890_),
    .A2(_02232_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10294_ (.A1(_03618_),
    .A2(_04630_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10295_ (.I(_04631_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10296_ (.I(_04589_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10297_ (.A1(_04076_),
    .A2(_04632_),
    .B1(_04633_),
    .B2(net191),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10298_ (.A1(_04632_),
    .A2(_04633_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10299_ (.A1(_03739_),
    .A2(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10300_ (.A1(_04629_),
    .A2(_04634_),
    .B1(_04636_),
    .B2(_01782_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10301_ (.A1(_04624_),
    .A2(_04637_),
    .B(_04401_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10302_ (.A1(_04624_),
    .A2(_04627_),
    .B(_04638_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10303_ (.A1(_04572_),
    .A2(_02956_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10304_ (.A1(_04572_),
    .A2(_04547_),
    .B(_04554_),
    .C(_04565_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10305_ (.A1(_04598_),
    .A2(_04639_),
    .B(_04603_),
    .C(_04621_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10306_ (.I(_04565_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10307_ (.A1(_03287_),
    .A2(_03291_),
    .A3(_03294_),
    .B1(_04575_),
    .B2(_03293_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10308_ (.I0(_03280_),
    .I1(_03281_),
    .S(_04643_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10309_ (.A1(_04572_),
    .A2(_04571_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10310_ (.A1(net202),
    .A2(_04589_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10311_ (.A1(_01793_),
    .A2(_04589_),
    .B(_04646_),
    .C(_04547_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10312_ (.A1(_04644_),
    .A2(_04645_),
    .B(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10313_ (.A1(_04124_),
    .A2(_04631_),
    .B1(_04569_),
    .B2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10314_ (.A1(_04642_),
    .A2(_04649_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10315_ (.A1(_01793_),
    .A2(_04640_),
    .B(_04641_),
    .C(_04650_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10316_ (.A1(_03652_),
    .A2(_02818_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10317_ (.A1(_01793_),
    .A2(_03653_),
    .B(_04623_),
    .C(_04652_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10318_ (.A1(_04545_),
    .A2(_04639_),
    .B1(_04651_),
    .B2(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10319_ (.A1(_04604_),
    .A2(_04620_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10320_ (.A1(_02205_),
    .A2(_04542_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10321_ (.A1(_02958_),
    .A2(_04655_),
    .B(_04644_),
    .C(_04656_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10322_ (.A1(_03613_),
    .A2(_04654_),
    .A3(_04657_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10323_ (.A1(_03127_),
    .A2(_04625_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10324_ (.A1(_01812_),
    .A2(_03749_),
    .B(_04658_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10325_ (.A1(_04172_),
    .A2(_04632_),
    .B1(_04633_),
    .B2(net206),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10326_ (.A1(_04580_),
    .A2(_04636_),
    .B1(_04660_),
    .B2(_04629_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10327_ (.A1(_04624_),
    .A2(_04661_),
    .B(_04401_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10328_ (.A1(_04624_),
    .A2(_04659_),
    .B(_04662_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10329_ (.I(_01513_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10330_ (.A1(_04218_),
    .A2(_04568_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10331_ (.A1(net207),
    .A2(_04633_),
    .B(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10332_ (.A1(_04663_),
    .A2(_04636_),
    .B1(_04665_),
    .B2(_04629_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10333_ (.A1(_04623_),
    .A2(_04666_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10334_ (.A1(_03752_),
    .A2(_04608_),
    .B(_04599_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10335_ (.A1(_01494_),
    .A2(_03753_),
    .B(_04622_),
    .C(_04668_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10336_ (.A1(_03613_),
    .A2(_04667_),
    .A3(_04669_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10337_ (.A1(_03235_),
    .A2(_03166_),
    .B(_03158_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10338_ (.A1(_03150_),
    .A2(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10339_ (.A1(_04656_),
    .A2(_04671_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10340_ (.A1(_01429_),
    .A2(_03665_),
    .Z(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10341_ (.A1(_01485_),
    .A2(_03585_),
    .B(_03368_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10342_ (.A1(_02816_),
    .A2(_04597_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10343_ (.A1(_01484_),
    .A2(_04588_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10344_ (.A1(_02333_),
    .A2(_04588_),
    .B(_04676_),
    .C(_03004_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10345_ (.A1(_01484_),
    .A2(_03298_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10346_ (.A1(_04580_),
    .A2(_01612_),
    .B(_02883_),
    .C(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10347_ (.A1(_02852_),
    .A2(_04677_),
    .A3(_04679_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10348_ (.A1(_04580_),
    .A2(_01642_),
    .B(_04678_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10349_ (.A1(_04581_),
    .A2(_04681_),
    .B(_04546_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10350_ (.A1(_04645_),
    .A2(_04671_),
    .B1(_04680_),
    .B2(_04682_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10351_ (.A1(_04259_),
    .A2(_04631_),
    .B1(_04569_),
    .B2(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(_04642_),
    .A2(_04684_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10353_ (.A1(_01485_),
    .A2(_04640_),
    .B(_04685_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10354_ (.I(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10355_ (.A1(_04656_),
    .A2(_04687_),
    .B(_04672_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10356_ (.A1(_04598_),
    .A2(_04674_),
    .B1(_04675_),
    .B2(_04688_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10357_ (.A1(_02816_),
    .A2(_04619_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10358_ (.A1(_01485_),
    .A2(_03756_),
    .A3(_04612_),
    .A4(_04690_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10359_ (.A1(_04689_),
    .A2(_04691_),
    .B(_04604_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10360_ (.A1(_04621_),
    .A2(_04620_),
    .A3(_04688_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10361_ (.A1(_04622_),
    .A2(_04687_),
    .A3(_04693_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10362_ (.A1(_04545_),
    .A2(_04639_),
    .B1(_04692_),
    .B2(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10363_ (.A1(_04672_),
    .A2(_04673_),
    .B(_04695_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10364_ (.A1(_03743_),
    .A2(_04696_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10365_ (.A1(_01458_),
    .A2(_02861_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10366_ (.A1(_04697_),
    .A2(_03273_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10367_ (.A1(_03137_),
    .A2(_03183_),
    .A3(_03231_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10368_ (.A1(_02892_),
    .A2(_02970_),
    .A3(_03031_),
    .A4(_03089_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10369_ (.A1(_04699_),
    .A2(_04700_),
    .ZN(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10370_ (.A1(_03662_),
    .A2(_03585_),
    .A3(_03655_),
    .A4(_03652_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10371_ (.A1(_03752_),
    .A2(_02973_),
    .A3(_04609_),
    .A4(_04702_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10372_ (.A1(_03761_),
    .A2(_04703_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10373_ (.I(_03728_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10374_ (.I(_02821_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10375_ (.A1(_02272_),
    .A2(_04706_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10376_ (.A1(_01861_),
    .A2(_04601_),
    .B(_02972_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10377_ (.I(_04600_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10378_ (.A1(net173),
    .A2(_04709_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10379_ (.A1(_01472_),
    .A2(_02954_),
    .B(_03265_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10380_ (.A1(_04707_),
    .A2(_04708_),
    .B1(_04710_),
    .B2(_04711_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10381_ (.A1(\as2650.debug_psu[5] ),
    .A2(_04709_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10382_ (.A1(_01484_),
    .A2(_02954_),
    .B(_03224_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10383_ (.A1(_02227_),
    .A2(_04706_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10384_ (.A1(_01851_),
    .A2(_01003_),
    .B(_02894_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10385_ (.A1(_04713_),
    .A2(_04714_),
    .B1(_04715_),
    .B2(_04716_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10386_ (.A1(\as2650.debug_psu[4] ),
    .A2(_04709_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10387_ (.A1(_01491_),
    .A2(_02954_),
    .B(_03172_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10388_ (.A1(_01811_),
    .A2(_04706_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10389_ (.A1(\as2650.debug_psu[3] ),
    .A2(_04601_),
    .B(_03127_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10390_ (.A1(_04718_),
    .A2(_04719_),
    .B1(_04720_),
    .B2(_04721_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10391_ (.A1(\as2650.debug_psl[7] ),
    .A2(_01001_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10392_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02820_),
    .B(_04723_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10393_ (.A1(\as2650.debug_psl[2] ),
    .A2(_04612_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10394_ (.A1(_01869_),
    .A2(_04601_),
    .B(_03080_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10395_ (.A1(_03275_),
    .A2(_04724_),
    .B1(_04725_),
    .B2(_04726_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10396_ (.A1(_04712_),
    .A2(_04717_),
    .A3(_04722_),
    .A4(_04727_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10397_ (.A1(_01428_),
    .A2(_03872_),
    .A3(_03624_),
    .Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10398_ (.A1(_04564_),
    .A2(_04548_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10399_ (.I(_04551_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10400_ (.A1(_02927_),
    .A2(_03001_),
    .A3(_03052_),
    .A4(_03112_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10401_ (.A1(_03166_),
    .A2(_03205_),
    .A3(_03249_),
    .A4(_04732_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10402_ (.A1(_04643_),
    .A2(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10403_ (.A1(_02834_),
    .A2(_01427_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10404_ (.A1(_02364_),
    .A2(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10405_ (.A1(_02348_),
    .A2(_02333_),
    .A3(_02316_),
    .A4(_01558_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10406_ (.A1(_01341_),
    .A2(_01349_),
    .A3(_01356_),
    .A4(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10407_ (.A1(_02815_),
    .A2(_01392_),
    .A3(_01397_),
    .A4(_02997_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10408_ (.I(net173),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10409_ (.A1(\as2650.debug_psu[5] ),
    .A2(\as2650.debug_psu[4] ),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10410_ (.A1(_02523_),
    .A2(_04740_),
    .A3(_02526_),
    .A4(_04741_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10411_ (.A1(_01506_),
    .A2(\as2650.debug_psl[6] ),
    .A3(\as2650.debug_psl[0] ),
    .A4(\as2650.debug_psl[5] ),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10412_ (.A1(_01782_),
    .A2(_01792_),
    .A3(_03298_),
    .A4(_04743_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10413_ (.A1(\as2650.debug_psu[7] ),
    .A2(_02819_),
    .A3(_04742_),
    .B1(_04744_),
    .B2(_04723_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10414_ (.A1(_00811_),
    .A2(_01397_),
    .A3(_01525_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10415_ (.I0(_04745_),
    .I1(_01471_),
    .S(_04746_),
    .Z(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10416_ (.A1(_01471_),
    .A2(_02819_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10417_ (.A1(_00637_),
    .A2(_02819_),
    .B(_04748_),
    .C(_04739_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10418_ (.A1(_04739_),
    .A2(_04747_),
    .B(_04749_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10419_ (.A1(_03207_),
    .A2(_03055_),
    .A3(_00932_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10420_ (.A1(_01050_),
    .A2(_02942_),
    .A3(_04751_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10421_ (.A1(_00984_),
    .A2(_02882_),
    .A3(_04752_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10422_ (.A1(_02882_),
    .A2(_04750_),
    .B(_04753_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10423_ (.A1(_02851_),
    .A2(_03301_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10424_ (.I(_00928_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10425_ (.A1(_04756_),
    .A2(_01567_),
    .A3(_01586_),
    .A4(_04751_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10426_ (.A1(_02852_),
    .A2(_04754_),
    .B1(_04755_),
    .B2(_04757_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10427_ (.A1(_04736_),
    .A2(_04738_),
    .B1(_04758_),
    .B2(_04735_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10428_ (.A1(_04570_),
    .A2(_04759_),
    .B(_04552_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10429_ (.A1(_04570_),
    .A2(_04734_),
    .B(_04760_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10430_ (.A1(_00633_),
    .A2(_04756_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10431_ (.A1(_01653_),
    .A2(_02941_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10432_ (.A1(_00642_),
    .A2(_01641_),
    .B(_04763_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10433_ (.A1(_00658_),
    .A2(_01611_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10434_ (.A1(_01632_),
    .A2(_03209_),
    .B(_04765_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10435_ (.A1(_01632_),
    .A2(_03209_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10436_ (.A1(_00658_),
    .A2(_01611_),
    .B1(_01356_),
    .B2(_01601_),
    .C(_04767_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10437_ (.A1(_04766_),
    .A2(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10438_ (.A1(_01586_),
    .A2(_01348_),
    .B1(_01356_),
    .B2(_01602_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10439_ (.A1(_01057_),
    .A2(_01331_),
    .B1(_01340_),
    .B2(_01567_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10440_ (.A1(_02936_),
    .A2(_02274_),
    .B(_04771_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10441_ (.A1(_01586_),
    .A2(_01348_),
    .B(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10442_ (.A1(_04770_),
    .A2(_04773_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _10443_ (.A1(_00642_),
    .A2(_01641_),
    .B1(_04766_),
    .B2(_04767_),
    .C1(_04769_),
    .C2(_04774_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10444_ (.A1(\as2650.debug_psl[1] ),
    .A2(_04763_),
    .B1(_04764_),
    .B2(_04775_),
    .C(_04762_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10445_ (.A1(_02271_),
    .A2(_04762_),
    .B(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _10446_ (.A1(net209),
    .A2(_01641_),
    .B1(_03299_),
    .B2(_01332_),
    .C1(_01341_),
    .C2(_01567_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10447_ (.A1(_01587_),
    .A2(_01349_),
    .B1(_01357_),
    .B2(_01602_),
    .C(_04771_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10448_ (.A1(_00633_),
    .A2(_04756_),
    .B1(_03059_),
    .B2(_01594_),
    .C(_04764_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10449_ (.A1(_04769_),
    .A2(_04778_),
    .A3(_04779_),
    .A4(_04780_),
    .Z(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10450_ (.A1(_04777_),
    .A2(_04781_),
    .B(_04553_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10451_ (.A1(_04731_),
    .A2(_04761_),
    .A3(_04782_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10452_ (.A1(_02464_),
    .A2(_02456_),
    .A3(_00645_),
    .A4(_01615_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10453_ (.A1(_00590_),
    .A2(_00649_),
    .B1(_00657_),
    .B2(_00585_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10454_ (.A1(_04784_),
    .A2(_04785_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10455_ (.A1(net184),
    .A2(_00640_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10456_ (.A1(_04786_),
    .A2(_04787_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10457_ (.A1(_04784_),
    .A2(_04788_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10458_ (.A1(net185),
    .A2(_00640_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10459_ (.A1(_00585_),
    .A2(_00649_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10460_ (.A1(_04790_),
    .A2(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10461_ (.A1(net184),
    .A2(_00631_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10462_ (.A1(_04792_),
    .A2(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10463_ (.A1(_04789_),
    .A2(_04794_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10464_ (.A1(_00584_),
    .A2(_01353_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10465_ (.A1(_00590_),
    .A2(_00656_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10466_ (.A1(_04797_),
    .A2(_04796_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _10467_ (.A1(_02456_),
    .A2(_01615_),
    .A3(_04796_),
    .B1(_04798_),
    .B2(_00645_),
    .B3(_02448_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10468_ (.A1(net183),
    .A2(_00632_),
    .B(net261),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10469_ (.A1(_04786_),
    .A2(_04787_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10470_ (.A1(net183),
    .A2(_00632_),
    .A3(net261),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10471_ (.A1(_04800_),
    .A2(_04801_),
    .B(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10472_ (.A1(_04795_),
    .A2(_04803_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10473_ (.A1(_04790_),
    .A2(_04791_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10474_ (.A1(_04792_),
    .A2(_04793_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10475_ (.A1(_00585_),
    .A2(_00641_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10476_ (.A1(net185),
    .A2(_00631_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10477_ (.A1(_04807_),
    .A2(_04808_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10478_ (.A1(_04805_),
    .A2(_04806_),
    .B(_04809_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10479_ (.A1(_04805_),
    .A2(_04806_),
    .A3(_04809_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10480_ (.A1(_04810_),
    .A2(_04811_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10481_ (.A1(_00602_),
    .A2(_00608_),
    .A3(_01329_),
    .A4(_01339_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10482_ (.I(_00600_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10483_ (.A1(_04814_),
    .A2(_01329_),
    .B1(_01338_),
    .B2(_00608_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10484_ (.I(_04815_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10485_ (.A1(_04813_),
    .A2(_04816_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10486_ (.A1(_00622_),
    .A2(_01353_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10487_ (.A1(_00614_),
    .A2(_01337_),
    .B1(_01346_),
    .B2(_00617_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10488_ (.I(_00611_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10489_ (.I(_04820_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10490_ (.A1(_04821_),
    .A2(_00617_),
    .A3(_01337_),
    .A4(_01346_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10491_ (.A1(_04818_),
    .A2(_04819_),
    .B(_04822_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10492_ (.A1(_00616_),
    .A2(_01351_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10493_ (.I(_01344_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10494_ (.A1(_04820_),
    .A2(_04825_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10495_ (.A1(_00622_),
    .A2(_00656_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10496_ (.A1(_04824_),
    .A2(_04826_),
    .A3(_04827_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10497_ (.A1(_04823_),
    .A2(_04828_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10498_ (.A1(_00614_),
    .A2(_00618_),
    .A3(_01328_),
    .A4(_01337_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10499_ (.A1(_00623_),
    .A2(_01346_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10500_ (.A1(_00614_),
    .A2(_01328_),
    .B1(_01338_),
    .B2(_00618_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10501_ (.A1(_04830_),
    .A2(_04831_),
    .A3(_04832_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10502_ (.A1(_00617_),
    .A2(_01345_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10503_ (.A1(_04821_),
    .A2(_01336_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10504_ (.A1(_04834_),
    .A2(_04835_),
    .A3(_04818_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10505_ (.A1(_04830_),
    .A2(_04833_),
    .B(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10506_ (.A1(_04829_),
    .A2(_04837_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10507_ (.A1(_04829_),
    .A2(_04837_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10508_ (.A1(_04817_),
    .A2(_04838_),
    .B(_04839_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10509_ (.A1(_02433_),
    .A2(_02421_),
    .A3(_02274_),
    .A4(_01343_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10510_ (.A1(_04814_),
    .A2(_01338_),
    .B1(_01348_),
    .B2(_00608_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10511_ (.A1(_04841_),
    .A2(_04842_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10512_ (.A1(_04823_),
    .A2(_04828_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10513_ (.I(_00615_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10514_ (.I(_04845_),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10515_ (.A1(_04821_),
    .A2(_04825_),
    .B1(_01352_),
    .B2(_04846_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10516_ (.A1(_04821_),
    .A2(_04846_),
    .A3(_04825_),
    .A4(_01352_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10517_ (.A1(_04827_),
    .A2(_04847_),
    .B(_04848_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10518_ (.A1(_00615_),
    .A2(_00654_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10519_ (.A1(_00612_),
    .A2(_01350_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10520_ (.A1(_00621_),
    .A2(_00647_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10521_ (.A1(_04850_),
    .A2(_04851_),
    .A3(_04852_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10522_ (.A1(_00596_),
    .A2(_01328_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10523_ (.A1(_04849_),
    .A2(_04853_),
    .A3(_04854_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10524_ (.A1(_04844_),
    .A2(_04855_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10525_ (.A1(_04843_),
    .A2(_04856_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10526_ (.A1(_04840_),
    .A2(_04857_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10527_ (.A1(_04813_),
    .A2(_04858_),
    .Z(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10528_ (.A1(_04830_),
    .A2(_04833_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10529_ (.A1(_04860_),
    .A2(_04836_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10530_ (.A1(_04830_),
    .A2(_04832_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10531_ (.A1(_04831_),
    .A2(_04862_),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10532_ (.A1(net212),
    .A2(_00623_),
    .A3(_01330_),
    .A4(_01339_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10533_ (.I(_04864_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10534_ (.A1(_04863_),
    .A2(_04865_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10535_ (.A1(_04861_),
    .A2(_04866_),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10536_ (.A1(_04861_),
    .A2(_04866_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10537_ (.A1(_00610_),
    .A2(_01330_),
    .A3(_04868_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10538_ (.A1(_04817_),
    .A2(_04838_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10539_ (.A1(_04867_),
    .A2(_04869_),
    .B(_04870_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10540_ (.A1(_04859_),
    .A2(_04871_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(_04840_),
    .A2(_04857_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10542_ (.A1(_04813_),
    .A2(_04858_),
    .B(_04873_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10543_ (.A1(_04844_),
    .A2(_04855_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10544_ (.A1(_04843_),
    .A2(_04856_),
    .B(_04875_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10545_ (.A1(_04849_),
    .A2(_04853_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10546_ (.A1(_04849_),
    .A2(_04853_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10547_ (.A1(_04854_),
    .A2(_04877_),
    .B(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10548_ (.A1(_00589_),
    .A2(_00594_),
    .A3(_01327_),
    .A4(_01336_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10549_ (.A1(_00589_),
    .A2(_01327_),
    .B1(_01336_),
    .B2(_00595_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10550_ (.A1(_04880_),
    .A2(_04881_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10551_ (.A1(_04845_),
    .A2(_00655_),
    .B1(_01351_),
    .B2(_00612_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10552_ (.A1(_04820_),
    .A2(_04845_),
    .A3(_00654_),
    .A4(_01350_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10553_ (.A1(_04852_),
    .A2(_04883_),
    .B(_04884_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10554_ (.A1(_00615_),
    .A2(_00646_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10555_ (.A1(_00611_),
    .A2(_00654_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10556_ (.A1(_00621_),
    .A2(_00638_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10557_ (.A1(_04886_),
    .A2(_04887_),
    .A3(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10558_ (.A1(_04885_),
    .A2(_04889_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10559_ (.A1(_04882_),
    .A2(_04890_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10560_ (.A1(_00600_),
    .A2(_00606_),
    .A3(_01347_),
    .A4(_01353_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10561_ (.A1(_00601_),
    .A2(_01347_),
    .B1(_01354_),
    .B2(_00607_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10562_ (.A1(_04892_),
    .A2(_04893_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10563_ (.A1(_04879_),
    .A2(_04891_),
    .A3(_04894_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10564_ (.A1(_04876_),
    .A2(_04895_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10565_ (.A1(_04841_),
    .A2(_04896_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10566_ (.A1(_04874_),
    .A2(_04897_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10567_ (.A1(_04874_),
    .A2(_04897_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10568_ (.A1(_04872_),
    .A2(_04898_),
    .B(_04899_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10569_ (.I(_04876_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10570_ (.A1(_04901_),
    .A2(_04895_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10571_ (.A1(_04841_),
    .A2(_04896_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10572_ (.A1(_04902_),
    .A2(_04903_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10573_ (.A1(_04879_),
    .A2(_04891_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10574_ (.A1(_04879_),
    .A2(_04891_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10575_ (.A1(_04892_),
    .A2(_04893_),
    .A3(_04905_),
    .B(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10576_ (.A1(_00607_),
    .A2(_00656_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10577_ (.A1(_00601_),
    .A2(_01354_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10578_ (.A1(_04880_),
    .A2(_04908_),
    .A3(_04909_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10579_ (.A1(_04885_),
    .A2(_04889_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10580_ (.A1(_04882_),
    .A2(_04890_),
    .B(_04911_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10581_ (.A1(_00595_),
    .A2(_01345_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10582_ (.A1(_00588_),
    .A2(_01335_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10583_ (.A1(_00583_),
    .A2(_01327_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10584_ (.A1(_04914_),
    .A2(_04915_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10585_ (.A1(_04913_),
    .A2(_04916_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10586_ (.A1(_00622_),
    .A2(_00629_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10587_ (.A1(_00612_),
    .A2(_04845_),
    .A3(_00638_),
    .A4(_00646_),
    .Z(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10588_ (.A1(_00616_),
    .A2(_00639_),
    .B1(_00647_),
    .B2(_04820_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10589_ (.A1(_04919_),
    .A2(_04920_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10590_ (.A1(_04846_),
    .A2(_00648_),
    .B1(_00655_),
    .B2(_00613_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10591_ (.A1(_00613_),
    .A2(_04846_),
    .A3(_00647_),
    .A4(_00655_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10592_ (.A1(_04888_),
    .A2(_04922_),
    .B(_04923_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10593_ (.A1(_04918_),
    .A2(_04921_),
    .A3(_04924_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10594_ (.A1(_04917_),
    .A2(_04925_),
    .Z(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10595_ (.A1(_04912_),
    .A2(_04926_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10596_ (.A1(_04910_),
    .A2(_04927_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10597_ (.A1(_04907_),
    .A2(_04928_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10598_ (.A1(_04892_),
    .A2(_04929_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10599_ (.A1(_04904_),
    .A2(_04930_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10600_ (.A1(_04904_),
    .A2(_04930_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10601_ (.A1(_04900_),
    .A2(_04931_),
    .B(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10602_ (.A1(_04907_),
    .A2(_04928_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10603_ (.A1(_04892_),
    .A2(_04929_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10604_ (.A1(_04934_),
    .A2(_04935_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10605_ (.A1(_00603_),
    .A2(_01355_),
    .B(_04880_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10606_ (.A1(_00603_),
    .A2(_01355_),
    .A3(_04880_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10607_ (.A1(_04908_),
    .A2(_04937_),
    .B(_04938_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10608_ (.A1(_04912_),
    .A2(_04926_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10609_ (.A1(_04910_),
    .A2(_04927_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10610_ (.A1(_04940_),
    .A2(_04941_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10611_ (.I(_04918_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10612_ (.A1(_04943_),
    .A2(_04921_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10613_ (.A1(_04924_),
    .A2(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10614_ (.A1(_04917_),
    .A2(_04925_),
    .B(_04945_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10615_ (.A1(_04943_),
    .A2(_04921_),
    .B(_04919_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10616_ (.A1(_00613_),
    .A2(_00639_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10617_ (.A1(_00616_),
    .A2(_00629_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10618_ (.A1(_04948_),
    .A2(_04949_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10619_ (.A1(_04948_),
    .A2(_04949_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10620_ (.A1(_04950_),
    .A2(_04951_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10621_ (.A1(_04947_),
    .A2(_04952_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10622_ (.A1(_00595_),
    .A2(_01352_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10623_ (.A1(_00588_),
    .A2(_04825_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10624_ (.A1(_00583_),
    .A2(_01335_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10625_ (.A1(_04955_),
    .A2(_04956_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10626_ (.A1(_04954_),
    .A2(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10627_ (.A1(_04953_),
    .A2(_04958_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10628_ (.A1(_04946_),
    .A2(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10629_ (.A1(_00609_),
    .A2(_00649_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10630_ (.A1(_00596_),
    .A2(_01347_),
    .A3(_04916_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10631_ (.A1(_04914_),
    .A2(_04915_),
    .B(_04962_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10632_ (.A1(_04814_),
    .A2(_00657_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10633_ (.A1(_04963_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10634_ (.A1(_04961_),
    .A2(_04965_),
    .Z(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10635_ (.A1(_04960_),
    .A2(_04966_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10636_ (.A1(_04942_),
    .A2(_04967_),
    .Z(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10637_ (.A1(_04939_),
    .A2(_04968_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10638_ (.A1(_04936_),
    .A2(_04969_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10639_ (.A1(_04936_),
    .A2(_04969_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10640_ (.A1(_04933_),
    .A2(_04970_),
    .B(_04971_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10641_ (.A1(_04942_),
    .A2(_04967_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10642_ (.A1(_04939_),
    .A2(_04968_),
    .B(_04973_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10643_ (.A1(_00602_),
    .A2(_00657_),
    .A3(_04963_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10644_ (.A1(_00610_),
    .A2(_00650_),
    .A3(_04965_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10645_ (.A1(_04975_),
    .A2(_04976_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10646_ (.A1(_04946_),
    .A2(_04959_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10647_ (.A1(_04960_),
    .A2(_04966_),
    .B(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10648_ (.A1(_04953_),
    .A2(_04958_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10649_ (.A1(_04947_),
    .A2(_04952_),
    .B(_04980_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10650_ (.A1(_02448_),
    .A2(_00653_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10651_ (.A1(_00589_),
    .A2(_01351_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10652_ (.A1(_00584_),
    .A2(_01345_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10653_ (.A1(_04982_),
    .A2(_04983_),
    .A3(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10654_ (.A1(_02393_),
    .A2(_00637_),
    .B(_00630_),
    .C(net181),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10655_ (.A1(_04985_),
    .A2(_04986_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10656_ (.A1(_04981_),
    .A2(_04987_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10657_ (.A1(_00609_),
    .A2(_00640_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10658_ (.A1(_02464_),
    .A2(_01334_),
    .A3(_04955_),
    .B1(_04957_),
    .B2(_04954_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10659_ (.A1(_00601_),
    .A2(_00648_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10660_ (.A1(_04990_),
    .A2(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10661_ (.A1(_04989_),
    .A2(_04992_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10662_ (.A1(_04988_),
    .A2(_04993_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10663_ (.A1(_04979_),
    .A2(_04994_),
    .Z(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10664_ (.A1(_04977_),
    .A2(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10665_ (.A1(_04974_),
    .A2(_04996_),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10666_ (.A1(_04974_),
    .A2(_04996_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10667_ (.A1(_04972_),
    .A2(_04997_),
    .B(_04998_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10668_ (.A1(_04979_),
    .A2(_04994_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10669_ (.A1(_04977_),
    .A2(_04995_),
    .B(_05000_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10670_ (.A1(_00603_),
    .A2(_00650_),
    .A3(_04990_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10671_ (.A1(_00610_),
    .A2(_00641_),
    .A3(_04992_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10672_ (.A1(_05002_),
    .A2(_05003_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10673_ (.A1(_04981_),
    .A2(_04987_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10674_ (.A1(_04988_),
    .A2(_04993_),
    .B(_05005_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10675_ (.A1(_04985_),
    .A2(_04986_),
    .B(_04950_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10676_ (.A1(_00596_),
    .A2(_00648_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10677_ (.A1(_04798_),
    .A2(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10678_ (.A1(_05007_),
    .A2(_05009_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10679_ (.A1(_00609_),
    .A2(_00630_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10680_ (.A1(_04983_),
    .A2(_04984_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10681_ (.A1(_04983_),
    .A2(_04984_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10682_ (.A1(_04982_),
    .A2(_05012_),
    .B(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10683_ (.A1(_04814_),
    .A2(_00639_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10684_ (.A1(_05014_),
    .A2(_05015_),
    .Z(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10685_ (.A1(_05011_),
    .A2(_05016_),
    .Z(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10686_ (.A1(_05010_),
    .A2(_05017_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10687_ (.A1(_05006_),
    .A2(_05018_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10688_ (.A1(_05004_),
    .A2(_05019_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10689_ (.A1(_05001_),
    .A2(_05020_),
    .Z(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10690_ (.I(_05001_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10691_ (.A1(_05022_),
    .A2(_05020_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10692_ (.A1(_04999_),
    .A2(_05021_),
    .B(_05023_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10693_ (.A1(_05006_),
    .A2(_05018_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10694_ (.A1(_05004_),
    .A2(_05019_),
    .B(_05025_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10695_ (.A1(net182),
    .A2(_00631_),
    .A3(_05016_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10696_ (.A1(_05014_),
    .A2(_05015_),
    .B(_05027_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10697_ (.I(_05009_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10698_ (.A1(_05010_),
    .A2(_05017_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10699_ (.A1(_05007_),
    .A2(_05029_),
    .B(_05030_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10700_ (.A1(_00602_),
    .A2(_00630_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10701_ (.A1(net262),
    .A2(_05032_),
    .A3(_04801_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10702_ (.A1(_05031_),
    .A2(_05033_),
    .Z(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10703_ (.A1(_05028_),
    .A2(_05034_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10704_ (.A1(_05026_),
    .A2(_05035_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10705_ (.A1(_05026_),
    .A2(_05035_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10706_ (.A1(_05024_),
    .A2(_05036_),
    .B(_05037_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10707_ (.A1(_05028_),
    .A2(_05034_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10708_ (.A1(_05031_),
    .A2(_05033_),
    .B(_05039_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10709_ (.A1(_04795_),
    .A2(_04803_),
    .Z(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10710_ (.A1(_05040_),
    .A2(_05041_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10711_ (.A1(_05040_),
    .A2(_05041_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10712_ (.A1(_05038_),
    .A2(_05042_),
    .B(_05043_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10713_ (.A1(_04789_),
    .A2(_04794_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10714_ (.I(_05045_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10715_ (.A1(_05046_),
    .A2(_04804_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10716_ (.A1(_04812_),
    .A2(_05047_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10717_ (.A1(_05044_),
    .A2(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10718_ (.A1(_04804_),
    .A2(_04812_),
    .B(_05049_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10719_ (.A1(net186),
    .A2(_00632_),
    .A3(_04790_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10720_ (.A1(_05046_),
    .A2(_04812_),
    .B(_04810_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10721_ (.A1(_05051_),
    .A2(_05052_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10722_ (.A1(_05050_),
    .A2(_05053_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10723_ (.A1(_05046_),
    .A2(_04812_),
    .B(_04810_),
    .C(_04790_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10724_ (.A1(net186),
    .A2(_00633_),
    .A3(_05055_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10725_ (.A1(_05054_),
    .A2(_05056_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10726_ (.A1(_04731_),
    .A2(_05057_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10727_ (.A1(_05050_),
    .A2(_05053_),
    .Z(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10728_ (.A1(_05044_),
    .A2(_05048_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10729_ (.A1(_05038_),
    .A2(_05042_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10730_ (.A1(_05024_),
    .A2(_05036_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10731_ (.A1(_04999_),
    .A2(_05021_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10732_ (.A1(_04972_),
    .A2(_04997_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _10733_ (.A1(_04936_),
    .A2(_04969_),
    .A3(_04933_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10734_ (.A1(_04900_),
    .A2(_04931_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10735_ (.A1(_04872_),
    .A2(_04898_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10736_ (.A1(_04859_),
    .A2(_04871_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10737_ (.A1(_04867_),
    .A2(_04869_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10738_ (.A1(_05069_),
    .A2(_04870_),
    .Z(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10739_ (.A1(net182),
    .A2(_01331_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10740_ (.A1(_05071_),
    .A2(_04868_),
    .Z(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10741_ (.A1(_04863_),
    .A2(_04864_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10742_ (.A1(net211),
    .A2(_01332_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10743_ (.A1(net212),
    .A2(_01331_),
    .B1(_01340_),
    .B2(_00623_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10744_ (.A1(_05072_),
    .A2(_05073_),
    .A3(_05074_),
    .A4(_05075_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10745_ (.A1(_05067_),
    .A2(_05068_),
    .A3(_05070_),
    .A4(_05076_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10746_ (.A1(_05064_),
    .A2(_05065_),
    .A3(_05066_),
    .A4(_05077_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10747_ (.A1(_05061_),
    .A2(_05062_),
    .A3(_05063_),
    .A4(_05078_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10748_ (.A1(_05059_),
    .A2(_05060_),
    .A3(_05079_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10749_ (.A1(_04549_),
    .A2(_04567_),
    .Z(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10750_ (.A1(_05058_),
    .A2(_05080_),
    .B(_05081_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10751_ (.A1(_04292_),
    .A2(_04567_),
    .B1(_04783_),
    .B2(_05082_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10752_ (.A1(_01471_),
    .A2(_04730_),
    .B1(_05083_),
    .B2(_04564_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10753_ (.A1(_02822_),
    .A2(_05084_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10754_ (.A1(_01472_),
    .A2(_03265_),
    .A3(_02822_),
    .Z(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10755_ (.A1(_05085_),
    .A2(_05086_),
    .B(_04690_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10756_ (.A1(_02164_),
    .A2(_03727_),
    .ZN(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _10757_ (.A1(_03655_),
    .A2(_01603_),
    .B1(_01587_),
    .B2(_03652_),
    .C1(_03366_),
    .C2(_03299_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10758_ (.A1(_03650_),
    .A2(_01568_),
    .B1(_01612_),
    .B2(_03144_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10759_ (.A1(_01678_),
    .A2(_03251_),
    .B1(_03208_),
    .B2(_03265_),
    .C(_05090_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10760_ (.A1(_03584_),
    .A2(_03138_),
    .B(_05091_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10761_ (.I(_02874_),
    .Z(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10762_ (.A1(_05088_),
    .A2(_05089_),
    .A3(_05092_),
    .B(_05093_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10763_ (.A1(_02875_),
    .A2(_05084_),
    .A3(_05094_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10764_ (.A1(_02955_),
    .A2(_04734_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10765_ (.A1(_05088_),
    .A2(_05096_),
    .B(_05094_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10766_ (.A1(_03274_),
    .A2(_01658_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10767_ (.A1(_03185_),
    .A2(_01636_),
    .B1(_01648_),
    .B2(_03489_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10768_ (.A1(_03457_),
    .A2(_01619_),
    .B1(_01636_),
    .B2(_03584_),
    .C(_05099_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10769_ (.A1(_03055_),
    .A2(_01652_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10770_ (.A1(_01652_),
    .A2(_01605_),
    .B(_05101_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10771_ (.I(_01619_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10772_ (.A1(_03127_),
    .A2(_05102_),
    .B1(_05103_),
    .B2(_03171_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(_01592_),
    .A2(_01595_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10774_ (.A1(_01587_),
    .A2(_01573_),
    .B(_05105_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10775_ (.A1(_03365_),
    .A2(_01561_),
    .B1(_01578_),
    .B2(_03401_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10776_ (.A1(_03650_),
    .A2(_01578_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10777_ (.A1(_03365_),
    .A2(_01561_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10778_ (.A1(_05108_),
    .A2(_05109_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10779_ (.A1(_03079_),
    .A2(_05106_),
    .B(_05107_),
    .C(_05110_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10780_ (.A1(_03079_),
    .A2(_05106_),
    .B1(_05102_),
    .B2(_03126_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10781_ (.A1(_03489_),
    .A2(_01648_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10782_ (.A1(_05112_),
    .A2(_05113_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10783_ (.A1(_05100_),
    .A2(_05104_),
    .A3(_05111_),
    .A4(_05114_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10784_ (.A1(_05098_),
    .A2(_05115_),
    .B(_05093_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10785_ (.A1(_03144_),
    .A2(_01619_),
    .B1(_01636_),
    .B2(_03584_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10786_ (.A1(_03079_),
    .A2(_05106_),
    .B1(_05107_),
    .B2(_05108_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10787_ (.A1(_05112_),
    .A2(_05118_),
    .B(_05104_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10788_ (.A1(_05117_),
    .A2(_05119_),
    .B(_05099_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10789_ (.A1(_05113_),
    .A2(_05120_),
    .B(_05098_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10790_ (.A1(_02271_),
    .A2(_03274_),
    .A3(_01658_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10791_ (.A1(_02271_),
    .A2(_03274_),
    .A3(_01658_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10792_ (.A1(_05121_),
    .A2(_05122_),
    .A3(_05123_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10793_ (.A1(_05116_),
    .A2(_05124_),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10794_ (.A1(_04675_),
    .A2(_05125_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10795_ (.A1(_01472_),
    .A2(_03662_),
    .B(_02822_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10796_ (.A1(_04606_),
    .A2(_05127_),
    .B(_04597_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10797_ (.A1(_05095_),
    .A2(_05097_),
    .A3(_05126_),
    .B1(_05128_),
    .B2(_05085_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10798_ (.A1(_05087_),
    .A2(_05129_),
    .ZN(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10799_ (.A1(_04705_),
    .A2(_05130_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10800_ (.A1(_04705_),
    .A2(_04728_),
    .B(_04729_),
    .C(_05131_),
    .ZN(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10801_ (.I(_04729_),
    .ZN(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10802_ (.I(_02957_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10803_ (.A1(_01429_),
    .A2(_05134_),
    .ZN(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10804_ (.A1(_05093_),
    .A2(_02956_),
    .B(_05135_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10805_ (.A1(_05084_),
    .A2(_05133_),
    .B(_05136_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10806_ (.A1(_05096_),
    .A2(_05125_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10807_ (.A1(_05132_),
    .A2(_05137_),
    .B1(_05138_),
    .B2(_04673_),
    .C(_02864_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10808_ (.A1(_02864_),
    .A2(_04704_),
    .B(_05139_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10809_ (.A1(_04698_),
    .A2(_04701_),
    .B1(_05140_),
    .B2(_04697_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10810_ (.A1(_03743_),
    .A2(_05141_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10811_ (.I(_05124_),
    .ZN(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10812_ (.A1(_04542_),
    .A2(_03296_),
    .B1(_05116_),
    .B2(_05142_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10813_ (.A1(_03630_),
    .A2(_03943_),
    .A3(_04642_),
    .ZN(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10814_ (.A1(_03296_),
    .A2(_04547_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10815_ (.A1(_02195_),
    .A2(_04586_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10816_ (.A1(\as2650.debug_psl[7] ),
    .A2(_04746_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10817_ (.A1(_04746_),
    .A2(_04724_),
    .B(_05147_),
    .C(_04739_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10818_ (.A1(net210),
    .A2(_04587_),
    .B1(_05146_),
    .B2(_01479_),
    .C(_05148_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10819_ (.A1(_03004_),
    .A2(_05149_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10820_ (.A1(_03208_),
    .A2(_03004_),
    .B(_05150_),
    .ZN(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10821_ (.A1(_02852_),
    .A2(_05151_),
    .B(_04755_),
    .ZN(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10822_ (.A1(_04735_),
    .A2(_05152_),
    .B(_04736_),
    .C(_04571_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10823_ (.A1(_05145_),
    .A2(_05153_),
    .B(_04553_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10824_ (.A1(_04553_),
    .A2(_04777_),
    .B(_05154_),
    .C(_04551_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _10825_ (.A1(_05081_),
    .A2(_05058_),
    .A3(_05155_),
    .B1(_04631_),
    .B2(_04338_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10826_ (.A1(_01479_),
    .A2(_05144_),
    .B1(_05156_),
    .B2(_04642_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10827_ (.A1(_05093_),
    .A2(_02956_),
    .A3(_04613_),
    .A4(_05088_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10828_ (.A1(_03761_),
    .A2(_04606_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10829_ (.A1(_01479_),
    .A2(_03761_),
    .B(_05159_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10830_ (.A1(_04613_),
    .A2(_05160_),
    .B(_05143_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10831_ (.A1(_04729_),
    .A2(_05161_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10832_ (.A1(_05157_),
    .A2(_05158_),
    .B(_05162_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10833_ (.A1(_04729_),
    .A2(_05157_),
    .ZN(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10834_ (.A1(_04705_),
    .A2(_05163_),
    .B(_05164_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10835_ (.A1(_05135_),
    .A2(_05143_),
    .B1(_05165_),
    .B2(_05136_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10836_ (.A1(_03075_),
    .A2(_05166_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10837_ (.A1(_03276_),
    .A2(_05167_),
    .B(_04698_),
    .C(_04275_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10838_ (.A1(_03771_),
    .A2(_03825_),
    .B(_02217_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10839_ (.A1(_04030_),
    .A2(_05168_),
    .B(_01852_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10840_ (.A1(_04706_),
    .A2(_04620_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10841_ (.I(_05170_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10842_ (.A1(_01852_),
    .A2(_04609_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10843_ (.A1(_04608_),
    .A2(_03736_),
    .B(_05172_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10844_ (.A1(_02217_),
    .A2(_03875_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10845_ (.A1(_05171_),
    .A2(_05173_),
    .B(_05174_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10846_ (.A1(_04621_),
    .A2(_05171_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10847_ (.I(_02261_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10848_ (.I(_04558_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10849_ (.A1(_05177_),
    .A2(_04313_),
    .A3(_05178_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10850_ (.I(_05146_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10851_ (.A1(_02251_),
    .A2(_05146_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10852_ (.A1(net180),
    .A2(_05180_),
    .B(_05181_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10853_ (.A1(_05179_),
    .A2(_05182_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10854_ (.A1(_03739_),
    .A2(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10855_ (.A1(_01852_),
    .A2(_03627_),
    .B(_05176_),
    .C(_05184_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10856_ (.A1(_02217_),
    .A2(_03769_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10857_ (.A1(_03764_),
    .A2(_05186_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10858_ (.A1(_01689_),
    .A2(_05175_),
    .B(_05185_),
    .C(_05187_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10859_ (.A1(_01463_),
    .A2(_05169_),
    .A3(_05188_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10860_ (.I(_05189_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10861_ (.I(_05187_),
    .Z(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10862_ (.A1(_02259_),
    .A2(_03906_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10863_ (.A1(_04602_),
    .A2(_01429_),
    .A3(_03624_),
    .A4(_04705_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10864_ (.A1(_01862_),
    .A2(_02973_),
    .B(_04626_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10865_ (.A1(_04599_),
    .A2(_05193_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10866_ (.A1(_02152_),
    .A2(_02218_),
    .A3(_05191_),
    .B1(_05192_),
    .B2(_05194_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10867_ (.A1(_04142_),
    .A2(_05195_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10868_ (.A1(_05171_),
    .A2(_05174_),
    .B(_03873_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10869_ (.A1(_04313_),
    .A2(_04558_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10870_ (.I(_03629_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10871_ (.A1(_02820_),
    .A2(_04739_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10872_ (.I(_05200_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10873_ (.I(_05200_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10874_ (.A1(net191),
    .A2(_05202_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10875_ (.A1(_02253_),
    .A2(_05201_),
    .B(_05203_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_02208_),
    .A2(_05199_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10877_ (.A1(_05199_),
    .A2(_05204_),
    .B1(_05205_),
    .B2(_01862_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10878_ (.A1(_05191_),
    .A2(_05198_),
    .B1(_05206_),
    .B2(_05178_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10879_ (.A1(_02478_),
    .A2(_05207_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10880_ (.A1(_05177_),
    .A2(_05191_),
    .B(_05208_),
    .C(_03627_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10881_ (.A1(_02253_),
    .A2(_03740_),
    .B(_05197_),
    .C(_05209_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10882_ (.A1(_05196_),
    .A2(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10883_ (.I(_01448_),
    .Z(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10884_ (.A1(_05191_),
    .A2(_05190_),
    .B(_05212_),
    .ZN(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10885_ (.A1(_05190_),
    .A2(_05211_),
    .B(_05213_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10886_ (.A1(_01868_),
    .A2(_02259_),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10887_ (.A1(_02218_),
    .A2(_05214_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10888_ (.A1(_02248_),
    .A2(_03653_),
    .B(_05170_),
    .C(_04652_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10889_ (.A1(_02152_),
    .A2(_05215_),
    .B(_05216_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10890_ (.A1(_05177_),
    .A2(_05214_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10891_ (.A1(net202),
    .A2(_05200_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10892_ (.A1(_02247_),
    .A2(_05202_),
    .B(_05219_),
    .ZN(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10893_ (.A1(_01869_),
    .A2(_05205_),
    .B1(_05220_),
    .B2(_05199_),
    .ZN(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10894_ (.A1(_03814_),
    .A2(_05198_),
    .B1(_05221_),
    .B2(_05178_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10895_ (.A1(_02478_),
    .A2(_05222_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10896_ (.A1(_05218_),
    .A2(_05223_),
    .B(_04628_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10897_ (.A1(_01871_),
    .A2(_03739_),
    .B(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10898_ (.A1(_04438_),
    .A2(_05217_),
    .B1(_05225_),
    .B2(_05197_),
    .C(_05186_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10899_ (.A1(_05186_),
    .A2(_05214_),
    .B(_05226_),
    .C(_03927_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10900_ (.A1(_03733_),
    .A2(_05215_),
    .B(_04401_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10901_ (.A1(_05227_),
    .A2(_05228_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10902_ (.A1(_01869_),
    .A2(_02259_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10903_ (.A1(_02615_),
    .A2(_05229_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10904_ (.A1(_01357_),
    .A2(_05202_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10905_ (.A1(_02523_),
    .A2(_05202_),
    .B(_05231_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10906_ (.A1(_01881_),
    .A2(_05205_),
    .B1(_05232_),
    .B2(_05199_),
    .ZN(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10907_ (.A1(_03782_),
    .A2(_05198_),
    .B1(_05233_),
    .B2(_05178_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10908_ (.A1(_02478_),
    .A2(_05234_),
    .Z(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10909_ (.A1(_05177_),
    .A2(_05230_),
    .B(_05235_),
    .C(_03616_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10910_ (.A1(_02524_),
    .A2(_04629_),
    .B(_05197_),
    .C(_05236_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10911_ (.A1(_01882_),
    .A2(_03128_),
    .B(_04658_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10912_ (.A1(_04599_),
    .A2(_05238_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10913_ (.A1(_02152_),
    .A2(_02218_),
    .A3(_05230_),
    .B1(_05239_),
    .B2(_05192_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10914_ (.A1(_04142_),
    .A2(_05240_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10915_ (.A1(_05237_),
    .A2(_05241_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10916_ (.A1(_05190_),
    .A2(_05230_),
    .B(_05212_),
    .ZN(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10917_ (.A1(_05190_),
    .A2(_05242_),
    .B(_05243_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10918_ (.I(_05176_),
    .Z(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10919_ (.I(_04568_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10920_ (.A1(_04524_),
    .A2(_05245_),
    .B1(_05201_),
    .B2(_02316_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10921_ (.A1(_04632_),
    .A2(_05180_),
    .B(_03711_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10922_ (.A1(_04352_),
    .A2(_05246_),
    .B1(_05247_),
    .B2(_01889_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10923_ (.A1(_01889_),
    .A2(_03752_),
    .B(_04668_),
    .C(_05192_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10924_ (.A1(_05244_),
    .A2(_05248_),
    .B1(_05249_),
    .B2(_04142_),
    .C(_01460_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _10925_ (.I(\as2650.debug_psu[5] ),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10926_ (.A1(_02215_),
    .A2(_04313_),
    .B1(_05180_),
    .B2(net208),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10927_ (.A1(_05250_),
    .A2(_05180_),
    .B1(_05251_),
    .B2(_04628_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10928_ (.A1(_04628_),
    .A2(_03822_),
    .A3(_04568_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10929_ (.A1(_01897_),
    .A2(_03616_),
    .B1(_05245_),
    .B2(_05252_),
    .C(_05253_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10930_ (.A1(_03660_),
    .A2(_02818_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10931_ (.A1(_05250_),
    .A2(_03660_),
    .B(_05171_),
    .C(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10932_ (.A1(_05244_),
    .A2(_05254_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10933_ (.A1(_01455_),
    .A2(_05256_),
    .B(_05257_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10934_ (.A1(_03608_),
    .A2(_05254_),
    .B(_05258_),
    .C(_03705_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10935_ (.A1(_03893_),
    .A2(_05245_),
    .B1(_05201_),
    .B2(_02348_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10936_ (.A1(_01903_),
    .A2(_05247_),
    .B1(_05259_),
    .B2(_04352_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10937_ (.A1(_03266_),
    .A2(_04608_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10938_ (.A1(_01903_),
    .A2(_03758_),
    .B(_05176_),
    .C(_05261_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10939_ (.A1(_05244_),
    .A2(_05260_),
    .B(_05262_),
    .C(_04275_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10940_ (.A1(_03921_),
    .A2(_05245_),
    .B1(_05201_),
    .B2(_02364_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10941_ (.A1(net37),
    .A2(_05247_),
    .B1(_05263_),
    .B2(_04352_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10942_ (.A1(_01910_),
    .A2(_03762_),
    .B(_05159_),
    .C(_05176_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10943_ (.I(_03963_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10944_ (.A1(_05244_),
    .A2(_05264_),
    .B(_05265_),
    .C(_05266_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10945_ (.A1(_03579_),
    .A2(_03700_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10946_ (.I(_05267_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10947_ (.I0(net44),
    .I1(\as2650.irqs_latch[1] ),
    .S(_05268_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10948_ (.I(_05269_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10949_ (.A1(net45),
    .A2(_05268_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10950_ (.A1(_01281_),
    .A2(_05268_),
    .B(_05270_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10951_ (.I0(net46),
    .I1(\as2650.irqs_latch[3] ),
    .S(_05268_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10952_ (.I(_05271_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10953_ (.I(_05267_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10954_ (.I0(\as2650.trap ),
    .I1(\as2650.irqs_latch[4] ),
    .S(_05272_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10955_ (.I(_05273_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10956_ (.I0(net47),
    .I1(\as2650.irqs_latch[5] ),
    .S(_05272_),
    .Z(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10957_ (.I(_05274_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10958_ (.I0(net48),
    .I1(\as2650.irqs_latch[6] ),
    .S(_05272_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10959_ (.I(_05275_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10960_ (.I0(net49),
    .I1(\as2650.irqs_latch[7] ),
    .S(_05272_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10961_ (.I(_05276_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10962_ (.A1(_03618_),
    .A2(_04555_),
    .A3(_04556_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10963_ (.A1(\as2650.trap ),
    .A2(_05277_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10964_ (.A1(_03618_),
    .A2(_04555_),
    .A3(_04550_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10965_ (.A1(_05278_),
    .A2(_05279_),
    .B(_03344_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10966_ (.I(_03717_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10967_ (.I(_05280_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10968_ (.I(_03718_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10969_ (.A1(net139),
    .A2(_05282_),
    .B(_05212_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10970_ (.A1(_03299_),
    .A2(_05281_),
    .B(_05283_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10971_ (.A1(net140),
    .A2(_05282_),
    .B(_05212_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10972_ (.A1(_01569_),
    .A2(_05281_),
    .B(_05284_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10973_ (.I(_03718_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10974_ (.I(_01448_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10975_ (.A1(net141),
    .A2(_05285_),
    .B(_05286_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10976_ (.A1(_01588_),
    .A2(_05281_),
    .B(_05287_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10977_ (.A1(net142),
    .A2(_05285_),
    .B(_05286_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10978_ (.A1(_01603_),
    .A2(_05281_),
    .B(_05288_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10979_ (.I(_05280_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10980_ (.A1(net143),
    .A2(_05285_),
    .B(_05286_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10981_ (.A1(_01613_),
    .A2(_05289_),
    .B(_05290_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10982_ (.A1(net144),
    .A2(_05285_),
    .B(_05286_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10983_ (.A1(_03138_),
    .A2(_05289_),
    .B(_05291_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10984_ (.A1(net145),
    .A2(_05280_),
    .B(_01449_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10985_ (.A1(_01642_),
    .A2(_05289_),
    .B(_05292_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10986_ (.A1(net146),
    .A2(_05280_),
    .B(_01449_),
    .ZN(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10987_ (.A1(_04756_),
    .A2(_05289_),
    .B(_05293_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10988_ (.A1(_00664_),
    .A2(_03693_),
    .B(net138),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10989_ (.A1(_03716_),
    .A2(_05282_),
    .A3(_05294_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10990_ (.I(_03730_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10991_ (.I(_05295_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10992_ (.A1(net132),
    .A2(_03731_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10993_ (.A1(_03736_),
    .A2(_05296_),
    .B(_05297_),
    .C(_05266_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10994_ (.A1(net133),
    .A2(_03731_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10995_ (.A1(_03744_),
    .A2(_05296_),
    .B(_05298_),
    .C(_05266_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10996_ (.A1(net134),
    .A2(_03731_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10997_ (.A1(_03081_),
    .A2(_05296_),
    .B(_05299_),
    .C(_05266_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10998_ (.I(_05295_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10999_ (.A1(net135),
    .A2(_05300_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11000_ (.I(_03519_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11001_ (.A1(_03749_),
    .A2(_05296_),
    .B(_05301_),
    .C(_05302_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11002_ (.I(_05295_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11003_ (.A1(net136),
    .A2(_05300_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11004_ (.A1(_03753_),
    .A2(_05303_),
    .B(_05304_),
    .C(_05302_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11005_ (.A1(net137),
    .A2(_05300_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11006_ (.A1(_03756_),
    .A2(_05303_),
    .B(_05305_),
    .C(_05302_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11007_ (.A1(_01438_),
    .A2(_05300_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11008_ (.A1(_03758_),
    .A2(_05303_),
    .B(_05306_),
    .C(_05302_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11009_ (.A1(_01437_),
    .A2(_05295_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11010_ (.A1(_03762_),
    .A2(_05303_),
    .B(_05307_),
    .C(_03613_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11011_ (.A1(\as2650.io_bus_we ),
    .A2(_03718_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11012_ (.A1(_01374_),
    .A2(_05282_),
    .B(_05308_),
    .C(_03716_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11013_ (.A1(_01531_),
    .A2(_00375_),
    .A3(_01541_),
    .Z(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11014_ (.I(_05309_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11015_ (.A1(_00713_),
    .A2(_01449_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11016_ (.A1(_03547_),
    .A2(_02201_),
    .A3(_03583_),
    .A4(_03368_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11017_ (.A1(_03356_),
    .A2(_02923_),
    .A3(_03548_),
    .A4(_05311_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11018_ (.A1(_02010_),
    .A2(_03580_),
    .B1(_05310_),
    .B2(_05312_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11019_ (.I(_01490_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11020_ (.A1(_05313_),
    .A2(_04625_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _11021_ (.A1(_04709_),
    .A2(_02886_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11022_ (.A1(_05314_),
    .A2(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11023_ (.I(_05316_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11024_ (.I(_02928_),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11025_ (.A1(_04602_),
    .A2(_02959_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11026_ (.A1(_05313_),
    .A2(_04625_),
    .A3(_05319_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11027_ (.I(_05320_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11028_ (.A1(_05314_),
    .A2(_05315_),
    .B(_05320_),
    .C(_02964_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11029_ (.I(_05322_),
    .Z(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11030_ (.A1(_05318_),
    .A2(_05321_),
    .B1(_05323_),
    .B2(\as2650.regs[2][0] ),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11031_ (.A1(_02953_),
    .A2(_05317_),
    .B(_05324_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11032_ (.I(_03002_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11033_ (.A1(_05325_),
    .A2(_05321_),
    .B1(_05323_),
    .B2(\as2650.regs[2][1] ),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11034_ (.A1(_03027_),
    .A2(_05317_),
    .B(_05326_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11035_ (.I(_03053_),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11036_ (.A1(_05327_),
    .A2(_05321_),
    .B1(_05323_),
    .B2(\as2650.regs[2][2] ),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11037_ (.A1(_03085_),
    .A2(_05317_),
    .B(_05328_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11038_ (.I(_03113_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11039_ (.A1(_05329_),
    .A2(_05321_),
    .B1(_05323_),
    .B2(\as2650.regs[2][3] ),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11040_ (.A1(_03132_),
    .A2(_05317_),
    .B(_05330_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11041_ (.I(_05316_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11042_ (.I(_03167_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11043_ (.I(_05320_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11044_ (.I(_05322_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11045_ (.A1(_05332_),
    .A2(_05333_),
    .B1(_05334_),
    .B2(\as2650.regs[2][4] ),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11046_ (.A1(_03178_),
    .A2(_05331_),
    .B(_05335_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11047_ (.I(_03206_),
    .Z(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11048_ (.A1(_05336_),
    .A2(_05333_),
    .B1(_05334_),
    .B2(\as2650.regs[2][5] ),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11049_ (.A1(_03228_),
    .A2(_05331_),
    .B(_05337_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11050_ (.I(_03250_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11051_ (.A1(_05338_),
    .A2(_05333_),
    .B1(_05334_),
    .B2(\as2650.regs[2][6] ),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11052_ (.A1(_03270_),
    .A2(_05331_),
    .B(_05339_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11053_ (.I(_03297_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11054_ (.A1(_05340_),
    .A2(_05333_),
    .B1(_05334_),
    .B2(\as2650.regs[2][7] ),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11055_ (.A1(_03316_),
    .A2(_05331_),
    .B(_05341_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11056_ (.I(_02232_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11057_ (.A1(_02230_),
    .A2(_02263_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11058_ (.I(_05343_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _11059_ (.A1(_01522_),
    .A2(_05342_),
    .A3(_05344_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11060_ (.A1(_04556_),
    .A2(_04630_),
    .B(_05344_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11061_ (.I(_05346_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11062_ (.A1(_02815_),
    .A2(_04600_),
    .A3(_05342_),
    .A4(_05343_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11063_ (.I(_05348_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11064_ (.A1(_02237_),
    .A2(_04560_),
    .A3(_04546_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11065_ (.I(_05350_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11066_ (.A1(_01527_),
    .A2(_02847_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11067_ (.I(_05352_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11068_ (.A1(_02237_),
    .A2(_04551_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11069_ (.I(_05354_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11070_ (.A1(_05351_),
    .A2(_05353_),
    .A3(_05355_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11071_ (.A1(_05345_),
    .A2(_05347_),
    .A3(_05349_),
    .A4(_05356_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11072_ (.A1(_01492_),
    .A2(_05357_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11073_ (.I(_05358_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11074_ (.A1(_02816_),
    .A2(_04600_),
    .A3(_05342_),
    .A4(_05344_),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11075_ (.I(_05360_),
    .Z(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11076_ (.I(_05361_),
    .Z(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11077_ (.I(_05345_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11078_ (.I(_05354_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11079_ (.I(_05352_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11080_ (.A1(_04630_),
    .A2(_05343_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11081_ (.I(_05366_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11082_ (.A1(net211),
    .A2(_05366_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11083_ (.I(_05352_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11084_ (.A1(_04013_),
    .A2(_05367_),
    .B(_05368_),
    .C(_05369_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11085_ (.A1(\as2650.chirpchar[0] ),
    .A2(_05365_),
    .B(_05355_),
    .C(_05370_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11086_ (.A1(_05074_),
    .A2(_05364_),
    .B(_05371_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11087_ (.I(_05350_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11088_ (.I0(_02928_),
    .I1(_05372_),
    .S(_05373_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11089_ (.A1(_05363_),
    .A2(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11090_ (.A1(_01522_),
    .A2(_05342_),
    .A3(_05344_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11091_ (.I(_05376_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11092_ (.I(_05360_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11093_ (.A1(_02228_),
    .A2(_05377_),
    .B(_05378_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11094_ (.A1(_02251_),
    .A2(_05362_),
    .B1(_05375_),
    .B2(_05379_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11095_ (.A1(_01513_),
    .A2(_01365_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11096_ (.A1(_01633_),
    .A2(_01652_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11097_ (.A1(_04542_),
    .A2(_05134_),
    .A3(_05381_),
    .A4(_05382_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11098_ (.A1(_02823_),
    .A2(_02824_),
    .A3(_02826_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11099_ (.A1(_02838_),
    .A2(_02849_),
    .A3(_03060_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11100_ (.A1(_03007_),
    .A2(_03015_),
    .A3(_03020_),
    .A4(_03006_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11101_ (.A1(_02866_),
    .A2(_05385_),
    .A3(_05386_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11102_ (.A1(_05384_),
    .A2(_05387_),
    .B(_04602_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11103_ (.A1(_02961_),
    .A2(_04607_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11104_ (.A1(_05388_),
    .A2(_05389_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11105_ (.I(_05390_),
    .Z(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11106_ (.A1(_05345_),
    .A2(_05347_),
    .A3(_05349_),
    .A4(_05356_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11107_ (.A1(_05313_),
    .A2(_05392_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11108_ (.I(_05393_),
    .Z(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11109_ (.A1(_01491_),
    .A2(_01366_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11110_ (.I(_05395_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11111_ (.I(_05396_),
    .Z(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11112_ (.A1(_01006_),
    .A2(_05397_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11113_ (.A1(_02951_),
    .A2(_05391_),
    .B(_05394_),
    .C(_05398_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11114_ (.A1(_05359_),
    .A2(_05380_),
    .B(_05383_),
    .C(_05399_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11115_ (.I(_05382_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11116_ (.A1(_04543_),
    .A2(_05134_),
    .A3(_05381_),
    .A4(_05401_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11117_ (.I(_05402_),
    .Z(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11118_ (.I(_05390_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11119_ (.I(_05381_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11120_ (.A1(_05393_),
    .A2(_05405_),
    .A3(_05383_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11121_ (.A1(_05404_),
    .A2(_05406_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11122_ (.I(_05407_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11123_ (.A1(_05318_),
    .A2(_05403_),
    .B1(_05408_),
    .B2(_00999_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11124_ (.A1(_05400_),
    .A2(_05409_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11125_ (.I(_05351_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11126_ (.A1(_02264_),
    .A2(_04731_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11127_ (.A1(_04864_),
    .A2(_05075_),
    .B(_05411_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11128_ (.I(_05366_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11129_ (.A1(_04076_),
    .A2(_05413_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11130_ (.A1(_02230_),
    .A2(_02264_),
    .A3(_04558_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11131_ (.I(_05415_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11132_ (.A1(net212),
    .A2(_05416_),
    .B(_05353_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11133_ (.A1(_01528_),
    .A2(_02847_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11134_ (.I(_05418_),
    .Z(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11135_ (.A1(\as2650.chirpchar[1] ),
    .A2(_05419_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11136_ (.I(_05354_),
    .Z(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11137_ (.A1(_05414_),
    .A2(_05417_),
    .B(_05420_),
    .C(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11138_ (.A1(_05412_),
    .A2(_05422_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11139_ (.A1(_05410_),
    .A2(_05423_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11140_ (.A1(_03002_),
    .A2(_05410_),
    .B(_05363_),
    .C(_05424_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11141_ (.A1(_02272_),
    .A2(_05377_),
    .B(_05378_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11142_ (.A1(_02253_),
    .A2(_05362_),
    .B1(_05425_),
    .B2(_05426_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11143_ (.A1(_01025_),
    .A2(_05397_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11144_ (.A1(_03025_),
    .A2(_05391_),
    .B(_05428_),
    .C(_05394_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11145_ (.I(_05383_),
    .Z(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11146_ (.A1(_05359_),
    .A2(_05427_),
    .B(_05429_),
    .C(_05430_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11147_ (.A1(_05325_),
    .A2(_05403_),
    .B1(_05408_),
    .B2(\as2650.regs[4][1] ),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11148_ (.A1(_05431_),
    .A2(_05432_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11149_ (.I(_05355_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11150_ (.A1(\as2650.chirpchar[2] ),
    .A2(_05419_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11151_ (.I(_05415_),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11152_ (.A1(_04124_),
    .A2(_05435_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11153_ (.A1(net181),
    .A2(_05435_),
    .B(_05436_),
    .C(_05369_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11154_ (.A1(_05434_),
    .A2(_05437_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11155_ (.A1(_05364_),
    .A2(_05438_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11156_ (.I(_05351_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11157_ (.A1(_05073_),
    .A2(_05433_),
    .B(_05439_),
    .C(_05440_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11158_ (.A1(_03053_),
    .A2(_05410_),
    .B(_05363_),
    .C(_05441_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11159_ (.A1(\as2650.debug_psl[2] ),
    .A2(_05376_),
    .B(_05361_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11160_ (.A1(_02249_),
    .A2(_05362_),
    .B1(_05442_),
    .B2(_05443_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11161_ (.I(_05390_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11162_ (.I(_05396_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11163_ (.A1(_01046_),
    .A2(_05446_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11164_ (.I(_05393_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11165_ (.A1(_03083_),
    .A2(_05445_),
    .B(_05447_),
    .C(_05448_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11166_ (.A1(_05359_),
    .A2(_05444_),
    .B(_05449_),
    .C(_05430_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11167_ (.A1(_05327_),
    .A2(_05403_),
    .B1(_05408_),
    .B2(\as2650.regs[4][2] ),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11168_ (.A1(_05450_),
    .A2(_05451_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11169_ (.I(_05345_),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11170_ (.A1(_04172_),
    .A2(_05367_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11171_ (.A1(net182),
    .A2(_05416_),
    .B(_05369_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11172_ (.A1(\as2650.chirpchar[3] ),
    .A2(_05418_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11173_ (.A1(_05453_),
    .A2(_05454_),
    .B(_05455_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11174_ (.A1(_05364_),
    .A2(_05456_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11175_ (.A1(_05072_),
    .A2(_05433_),
    .B(_05457_),
    .C(_05440_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11176_ (.A1(_03113_),
    .A2(_05410_),
    .B(_05452_),
    .C(_05458_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11177_ (.A1(_01812_),
    .A2(_05376_),
    .B(_05361_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11178_ (.A1(_02524_),
    .A2(_05362_),
    .B1(_05459_),
    .B2(_05460_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11179_ (.A1(\as2650.regs[0][3] ),
    .A2(_05446_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11180_ (.A1(_03130_),
    .A2(_05445_),
    .B(_05462_),
    .C(_05448_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11181_ (.A1(_05359_),
    .A2(_05461_),
    .B(_05463_),
    .C(_05430_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11182_ (.I(_05402_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11183_ (.I(_05407_),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11184_ (.A1(_05329_),
    .A2(_05465_),
    .B1(_05466_),
    .B2(\as2650.regs[4][3] ),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11185_ (.A1(_05464_),
    .A2(_05467_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11186_ (.I(_05361_),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11187_ (.A1(_01889_),
    .A2(_05468_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11188_ (.I(_05452_),
    .Z(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11189_ (.I(_05373_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11190_ (.I(_05421_),
    .Z(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11191_ (.A1(net183),
    .A2(_05367_),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11192_ (.A1(_04218_),
    .A2(_05413_),
    .B(_05473_),
    .C(_05353_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11193_ (.A1(\as2650.chirpchar[4] ),
    .A2(_05365_),
    .B(_05364_),
    .C(_05474_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11194_ (.A1(_05070_),
    .A2(_05472_),
    .B(_05475_),
    .C(_05440_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11195_ (.A1(_03167_),
    .A2(_05471_),
    .B(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11196_ (.A1(_05470_),
    .A2(_05477_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11197_ (.A1(_01493_),
    .A2(_05470_),
    .B(_05349_),
    .C(_05478_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11198_ (.A1(_05469_),
    .A2(_05479_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11199_ (.A1(\as2650.regs[0][4] ),
    .A2(_05446_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11200_ (.A1(_03177_),
    .A2(_05445_),
    .B(_05481_),
    .C(_05448_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11201_ (.A1(_05358_),
    .A2(_05480_),
    .B(_05482_),
    .C(_05430_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11202_ (.A1(_05332_),
    .A2(_05465_),
    .B1(_05466_),
    .B2(\as2650.regs[4][4] ),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11203_ (.A1(_05483_),
    .A2(_05484_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11204_ (.I(_05421_),
    .Z(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11205_ (.A1(_04259_),
    .A2(_05413_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11206_ (.I(_05435_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11207_ (.A1(net184),
    .A2(_05487_),
    .B(_05365_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11208_ (.A1(\as2650.chirpchar[5] ),
    .A2(_05419_),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11209_ (.A1(_05486_),
    .A2(_05488_),
    .B(_05489_),
    .ZN(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11210_ (.A1(_05485_),
    .A2(_05490_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11211_ (.A1(_05068_),
    .A2(_05485_),
    .B(_05491_),
    .C(_05471_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11212_ (.A1(_03206_),
    .A2(_05471_),
    .B(_05470_),
    .C(_05492_),
    .ZN(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11213_ (.A1(_01486_),
    .A2(_05377_),
    .B(_05468_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _11214_ (.A1(_05250_),
    .A2(_05468_),
    .B1(_05493_),
    .B2(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11215_ (.A1(\as2650.regs[0][5] ),
    .A2(_05446_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11216_ (.A1(_03227_),
    .A2(_05445_),
    .B(_05496_),
    .C(_05448_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11217_ (.A1(_05358_),
    .A2(_05495_),
    .B(_05497_),
    .C(_05383_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11218_ (.A1(_05336_),
    .A2(_05465_),
    .B1(_05466_),
    .B2(\as2650.regs[4][5] ),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11219_ (.A1(_05498_),
    .A2(_05499_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11220_ (.A1(\as2650.regs[4][6] ),
    .A2(_05408_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11221_ (.A1(_04544_),
    .A2(_04545_),
    .A3(_05405_),
    .A4(_05401_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11222_ (.A1(\as2650.regs[0][6] ),
    .A2(_05397_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11223_ (.A1(_03269_),
    .A2(_05391_),
    .B(_05502_),
    .C(_05394_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11224_ (.A1(_04291_),
    .A2(_05367_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11225_ (.A1(net185),
    .A2(_05416_),
    .B(_05353_),
    .ZN(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11226_ (.A1(\as2650.chirpchar[6] ),
    .A2(_05419_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11227_ (.A1(_05504_),
    .A2(_05505_),
    .B(_05506_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11228_ (.A1(_05433_),
    .A2(_05507_),
    .ZN(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11229_ (.A1(_05067_),
    .A2(_05472_),
    .B(_05508_),
    .C(_05440_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11230_ (.A1(_03250_),
    .A2(_05471_),
    .B(_05363_),
    .C(_05509_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11231_ (.A1(_01473_),
    .A2(_05377_),
    .B(_05378_),
    .ZN(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _11232_ (.A1(_04740_),
    .A2(_05468_),
    .B1(_05510_),
    .B2(_05511_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11233_ (.A1(_05393_),
    .A2(_05512_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11234_ (.A1(_05501_),
    .A2(_05513_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11235_ (.A1(_05338_),
    .A2(_05501_),
    .B1(_05503_),
    .B2(_05514_),
    .ZN(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11236_ (.A1(_05500_),
    .A2(_05515_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11237_ (.I(_05394_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11238_ (.A1(net186),
    .A2(_05435_),
    .B(_05355_),
    .C(_05369_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11239_ (.A1(_04338_),
    .A2(_05416_),
    .B(_05517_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11240_ (.A1(_05066_),
    .A2(_05411_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11241_ (.A1(_05351_),
    .A2(_05519_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11242_ (.A1(_03297_),
    .A2(_05373_),
    .B1(_05518_),
    .B2(_05520_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11243_ (.A1(_05452_),
    .A2(_05521_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11244_ (.A1(_01480_),
    .A2(_05470_),
    .B(_05349_),
    .C(_05522_),
    .ZN(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11245_ (.A1(_01910_),
    .A2(_05378_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11246_ (.A1(_05523_),
    .A2(_05524_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11247_ (.A1(\as2650.regs[0][7] ),
    .A2(_05397_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11248_ (.A1(_03314_),
    .A2(_05391_),
    .B(_05526_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11249_ (.A1(_05516_),
    .A2(_05525_),
    .B(_05527_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11250_ (.A1(_05340_),
    .A2(_05465_),
    .B1(_05466_),
    .B2(\as2650.regs[4][7] ),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11251_ (.A1(_05403_),
    .A2(_05528_),
    .B(_05529_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11252_ (.A1(_01513_),
    .A2(_02886_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11253_ (.A1(_00890_),
    .A2(_05530_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11254_ (.I(_05531_),
    .Z(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11255_ (.A1(_01491_),
    .A2(_02817_),
    .A3(_02960_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11256_ (.I(_05533_),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11257_ (.I(_05411_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11258_ (.I(_05535_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11259_ (.A1(_05065_),
    .A2(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11260_ (.I(_05487_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11261_ (.I(_05538_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11262_ (.I(_05487_),
    .Z(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11263_ (.A1(_04388_),
    .A2(_05540_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11264_ (.I(_05485_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11265_ (.A1(net180),
    .A2(_05539_),
    .B(_05541_),
    .C(_05542_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11266_ (.A1(_05537_),
    .A2(_05543_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11267_ (.A1(_05433_),
    .A2(_05347_),
    .B(_02961_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11268_ (.I(_05545_),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11269_ (.A1(_01367_),
    .A2(_05545_),
    .A3(_05533_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11270_ (.A1(_05547_),
    .A2(_05531_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11271_ (.I(_05548_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11272_ (.A1(_02967_),
    .A2(_05534_),
    .B1(_05544_),
    .B2(_05546_),
    .C1(_05549_),
    .C2(\as2650.regs[1][0] ),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11273_ (.A1(_02953_),
    .A2(_05532_),
    .B(_05550_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11274_ (.A1(_05064_),
    .A2(_05536_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11275_ (.I(_05487_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11276_ (.A1(_04426_),
    .A2(_05552_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11277_ (.A1(net191),
    .A2(_05539_),
    .B(_05553_),
    .C(_05542_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11278_ (.A1(_05551_),
    .A2(_05554_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11279_ (.A1(_03028_),
    .A2(_05534_),
    .B1(_05555_),
    .B2(_05546_),
    .C1(_05549_),
    .C2(\as2650.regs[1][1] ),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11280_ (.A1(_03027_),
    .A2(_05532_),
    .B(_05556_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11281_ (.A1(_04445_),
    .A2(_04452_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11282_ (.A1(_05557_),
    .A2(_05538_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11283_ (.A1(net202),
    .A2(_05413_),
    .B(_05558_),
    .C(_05535_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11284_ (.A1(_05063_),
    .A2(_05536_),
    .B(_05559_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11285_ (.A1(_03086_),
    .A2(_05534_),
    .B1(_05560_),
    .B2(_05546_),
    .C1(_05549_),
    .C2(\as2650.regs[1][2] ),
    .ZN(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11286_ (.A1(_03085_),
    .A2(_05532_),
    .B(_05561_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11287_ (.A1(_04487_),
    .A2(_05538_),
    .ZN(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11288_ (.I(_05472_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11289_ (.A1(net206),
    .A2(_05540_),
    .B(_05562_),
    .C(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _11290_ (.A1(_05062_),
    .A2(_05542_),
    .B(_05564_),
    .ZN(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11291_ (.A1(_03133_),
    .A2(_05534_),
    .B1(_05565_),
    .B2(_05546_),
    .C1(_05549_),
    .C2(\as2650.regs[1][3] ),
    .ZN(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11292_ (.A1(_03132_),
    .A2(_05532_),
    .B(_05566_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11293_ (.I(_05531_),
    .Z(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11294_ (.I(_05533_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11295_ (.A1(_04524_),
    .A2(_05538_),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11296_ (.A1(net207),
    .A2(_05540_),
    .B(_05569_),
    .C(_05485_),
    .ZN(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _11297_ (.A1(_05061_),
    .A2(_05542_),
    .B(_05570_),
    .ZN(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11298_ (.I(_05545_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11299_ (.I(_05548_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11300_ (.A1(_03180_),
    .A2(_05568_),
    .B1(_05571_),
    .B2(_05572_),
    .C1(_05573_),
    .C2(\as2650.regs[1][4] ),
    .ZN(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11301_ (.A1(_03178_),
    .A2(_05567_),
    .B(_05574_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11302_ (.A1(_05060_),
    .A2(_05536_),
    .ZN(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11303_ (.A1(_03822_),
    .A2(_05552_),
    .ZN(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11304_ (.A1(net208),
    .A2(_05539_),
    .B(_05576_),
    .C(_05563_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11305_ (.A1(_05575_),
    .A2(_05577_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11306_ (.A1(_03229_),
    .A2(_05568_),
    .B1(_05578_),
    .B2(_05572_),
    .C1(_05573_),
    .C2(\as2650.regs[1][5] ),
    .ZN(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11307_ (.A1(_03228_),
    .A2(_05567_),
    .B(_05579_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11308_ (.A1(_05059_),
    .A2(_05535_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11309_ (.A1(_03893_),
    .A2(_05552_),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11310_ (.A1(net209),
    .A2(_05539_),
    .B(_05581_),
    .C(_05563_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11311_ (.A1(_05580_),
    .A2(_05582_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11312_ (.A1(_03271_),
    .A2(_05568_),
    .B1(_05583_),
    .B2(_05572_),
    .C1(_05573_),
    .C2(\as2650.regs[1][6] ),
    .ZN(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11313_ (.A1(_03270_),
    .A2(_05567_),
    .B(_05584_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11314_ (.A1(_05057_),
    .A2(_05535_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11315_ (.A1(_03921_),
    .A2(_05552_),
    .ZN(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11316_ (.A1(net210),
    .A2(_05540_),
    .B(_05586_),
    .C(_05563_),
    .ZN(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11317_ (.A1(_05585_),
    .A2(_05587_),
    .ZN(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11318_ (.A1(_03317_),
    .A2(_05568_),
    .B1(_05588_),
    .B2(_05572_),
    .C1(_05573_),
    .C2(\as2650.regs[1][7] ),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11319_ (.A1(_03316_),
    .A2(_05567_),
    .B(_05589_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11320_ (.A1(_03368_),
    .A2(_05530_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11321_ (.I(_05590_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11322_ (.A1(_02961_),
    .A2(_04607_),
    .A3(_02960_),
    .ZN(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11323_ (.I(_05592_),
    .Z(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11324_ (.A1(_02964_),
    .A2(_05592_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11325_ (.A1(_05594_),
    .A2(_05590_),
    .Z(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11326_ (.I(_05595_),
    .Z(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11327_ (.A1(_05318_),
    .A2(_05593_),
    .B1(_05596_),
    .B2(\as2650.regs[3][0] ),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11328_ (.A1(_02953_),
    .A2(_05591_),
    .B(_05597_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11329_ (.A1(_05325_),
    .A2(_05593_),
    .B1(_05596_),
    .B2(\as2650.regs[3][1] ),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11330_ (.A1(_03027_),
    .A2(_05591_),
    .B(_05598_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11331_ (.A1(_05327_),
    .A2(_05593_),
    .B1(_05596_),
    .B2(\as2650.regs[3][2] ),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11332_ (.A1(_03085_),
    .A2(_05591_),
    .B(_05599_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11333_ (.A1(_05329_),
    .A2(_05593_),
    .B1(_05596_),
    .B2(\as2650.regs[3][3] ),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11334_ (.A1(_03132_),
    .A2(_05591_),
    .B(_05600_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11335_ (.I(_05590_),
    .Z(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11336_ (.I(_05592_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11337_ (.I(_05595_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11338_ (.A1(_05332_),
    .A2(_05602_),
    .B1(_05603_),
    .B2(\as2650.regs[3][4] ),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11339_ (.A1(_03178_),
    .A2(_05601_),
    .B(_05604_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11340_ (.A1(_05336_),
    .A2(_05602_),
    .B1(_05603_),
    .B2(\as2650.regs[3][5] ),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11341_ (.A1(_03228_),
    .A2(_05601_),
    .B(_05605_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11342_ (.A1(_05338_),
    .A2(_05602_),
    .B1(_05603_),
    .B2(\as2650.regs[3][6] ),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11343_ (.A1(_03270_),
    .A2(_05601_),
    .B(_05606_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11344_ (.A1(_05340_),
    .A2(_05602_),
    .B1(_05603_),
    .B2(\as2650.regs[3][7] ),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11345_ (.A1(_03316_),
    .A2(_05601_),
    .B(_05607_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11346_ (.A1(_04607_),
    .A2(_02887_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11347_ (.I(_05608_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11348_ (.A1(_05472_),
    .A2(_05347_),
    .B(_04663_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11349_ (.I(_05610_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11350_ (.A1(_02960_),
    .A2(_05389_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11351_ (.I(_05612_),
    .Z(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11352_ (.I(_05608_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _11353_ (.A1(_02964_),
    .A2(_05610_),
    .A3(_05612_),
    .A4(_05614_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11354_ (.I(_05615_),
    .Z(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11355_ (.A1(_05544_),
    .A2(_05611_),
    .B1(_05613_),
    .B2(_02967_),
    .C1(\as2650.regs[5][0] ),
    .C2(_05616_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11356_ (.A1(_02952_),
    .A2(_05609_),
    .B(_05617_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11357_ (.A1(_05555_),
    .A2(_05611_),
    .B1(_05613_),
    .B2(_03028_),
    .C1(\as2650.regs[5][1] ),
    .C2(_05616_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11358_ (.A1(_03026_),
    .A2(_05609_),
    .B(_05618_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11359_ (.A1(_05560_),
    .A2(_05611_),
    .B1(_05613_),
    .B2(_03086_),
    .C1(\as2650.regs[5][2] ),
    .C2(_05616_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11360_ (.A1(_03084_),
    .A2(_05609_),
    .B(_05619_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11361_ (.A1(_05565_),
    .A2(_05611_),
    .B1(_05613_),
    .B2(_03133_),
    .C1(\as2650.regs[5][3] ),
    .C2(_05616_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11362_ (.A1(_03131_),
    .A2(_05609_),
    .B(_05620_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11363_ (.I(_05608_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11364_ (.I(_05610_),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11365_ (.I(_05612_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11366_ (.I(_05615_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11367_ (.A1(_05571_),
    .A2(_05622_),
    .B1(_05623_),
    .B2(_03180_),
    .C1(\as2650.regs[5][4] ),
    .C2(_05624_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11368_ (.A1(_03177_),
    .A2(_05621_),
    .B(_05625_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11369_ (.A1(_05578_),
    .A2(_05622_),
    .B1(_05623_),
    .B2(_03229_),
    .C1(\as2650.regs[5][5] ),
    .C2(_05624_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11370_ (.A1(_03227_),
    .A2(_05621_),
    .B(_05626_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11371_ (.A1(_05583_),
    .A2(_05622_),
    .B1(_05623_),
    .B2(_03271_),
    .C1(\as2650.regs[5][6] ),
    .C2(_05624_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11372_ (.A1(_03269_),
    .A2(_05621_),
    .B(_05627_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11373_ (.A1(_05588_),
    .A2(_05622_),
    .B1(_05623_),
    .B2(_03317_),
    .C1(\as2650.regs[5][7] ),
    .C2(_05624_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11374_ (.A1(_03315_),
    .A2(_05621_),
    .B(_05628_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11375_ (.A1(_05313_),
    .A2(_02817_),
    .A3(_05315_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11376_ (.I(_05629_),
    .Z(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11377_ (.A1(_02962_),
    .A2(_05319_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11378_ (.I(_05631_),
    .Z(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11379_ (.I(_05629_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11380_ (.A1(_03518_),
    .A2(_05631_),
    .A3(_05633_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11381_ (.I(_05634_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11382_ (.A1(_02967_),
    .A2(_05632_),
    .B1(_05635_),
    .B2(\as2650.regs[6][0] ),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11383_ (.A1(_02952_),
    .A2(_05630_),
    .B(_05636_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11384_ (.A1(_03028_),
    .A2(_05632_),
    .B1(_05635_),
    .B2(\as2650.regs[6][1] ),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11385_ (.A1(_03026_),
    .A2(_05630_),
    .B(_05637_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11386_ (.A1(_03086_),
    .A2(_05632_),
    .B1(_05635_),
    .B2(\as2650.regs[6][2] ),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11387_ (.A1(_03084_),
    .A2(_05630_),
    .B(_05638_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11388_ (.A1(_03133_),
    .A2(_05632_),
    .B1(_05635_),
    .B2(\as2650.regs[6][3] ),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11389_ (.A1(_03131_),
    .A2(_05630_),
    .B(_05639_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11390_ (.I(_05629_),
    .Z(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11391_ (.I(_05631_),
    .Z(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11392_ (.I(_05634_),
    .Z(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11393_ (.A1(_03180_),
    .A2(_05641_),
    .B1(_05642_),
    .B2(\as2650.regs[6][4] ),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11394_ (.A1(_03177_),
    .A2(_05640_),
    .B(_05643_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11395_ (.A1(_03229_),
    .A2(_05641_),
    .B1(_05642_),
    .B2(\as2650.regs[6][5] ),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11396_ (.A1(_03227_),
    .A2(_05640_),
    .B(_05644_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11397_ (.A1(_03271_),
    .A2(_05641_),
    .B1(_05642_),
    .B2(\as2650.regs[6][6] ),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11398_ (.A1(_03269_),
    .A2(_05640_),
    .B(_05645_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11399_ (.A1(_03317_),
    .A2(_05641_),
    .B1(_05642_),
    .B2(\as2650.regs[6][7] ),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11400_ (.A1(_03315_),
    .A2(_05640_),
    .B(_05646_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11401_ (.A1(_04543_),
    .A2(_05134_),
    .A3(_05395_),
    .A4(_05401_),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11402_ (.I(_05647_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11403_ (.A1(_02231_),
    .A2(_05530_),
    .ZN(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11404_ (.I(_05649_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11405_ (.I(_05405_),
    .Z(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11406_ (.A1(_05365_),
    .A2(_05421_),
    .A3(_05346_),
    .A4(_05348_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11407_ (.A1(_05373_),
    .A2(_05452_),
    .A3(_05652_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11408_ (.A1(_04663_),
    .A2(_05653_),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11409_ (.I(_05654_),
    .Z(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11410_ (.A1(_00999_),
    .A2(_05651_),
    .B1(_05380_),
    .B2(_05655_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11411_ (.A1(_02952_),
    .A2(_05650_),
    .B(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11412_ (.A1(_05648_),
    .A2(_05657_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _11413_ (.A1(_04543_),
    .A2(_03665_),
    .A3(_05396_),
    .A4(_05401_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11414_ (.I(_05659_),
    .Z(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11415_ (.A1(_04663_),
    .A2(_05357_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11416_ (.A1(_05396_),
    .A2(_05647_),
    .A3(_05661_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11417_ (.A1(_02231_),
    .A2(_05530_),
    .B(_05662_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11418_ (.I(_05663_),
    .Z(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11419_ (.A1(_05318_),
    .A2(_05660_),
    .B1(_05664_),
    .B2(_01006_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11420_ (.A1(_05658_),
    .A2(_05665_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11421_ (.A1(\as2650.regs[4][1] ),
    .A2(_05651_),
    .B1(_05427_),
    .B2(_05655_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11422_ (.A1(_03026_),
    .A2(_05650_),
    .B(_05666_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11423_ (.A1(_05648_),
    .A2(_05667_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11424_ (.A1(_05325_),
    .A2(_05660_),
    .B1(_05664_),
    .B2(_01025_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11425_ (.A1(_05668_),
    .A2(_05669_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11426_ (.A1(\as2650.regs[4][2] ),
    .A2(_05651_),
    .B1(_05444_),
    .B2(_05655_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11427_ (.A1(_03084_),
    .A2(_05650_),
    .B(_05670_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11428_ (.A1(_05648_),
    .A2(_05671_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11429_ (.A1(_05327_),
    .A2(_05660_),
    .B1(_05664_),
    .B2(_01046_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11430_ (.A1(_05672_),
    .A2(_05673_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11431_ (.A1(\as2650.regs[4][3] ),
    .A2(_05651_),
    .B1(_05461_),
    .B2(_05655_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11432_ (.A1(_03131_),
    .A2(_05650_),
    .B(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11433_ (.A1(_05648_),
    .A2(_05675_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11434_ (.A1(_05329_),
    .A2(_05660_),
    .B1(_05664_),
    .B2(\as2650.regs[0][3] ),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11435_ (.A1(_05676_),
    .A2(_05677_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11436_ (.I(_05661_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11437_ (.I(_05649_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11438_ (.I(_05405_),
    .Z(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11439_ (.A1(\as2650.regs[4][4] ),
    .A2(_05680_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11440_ (.A1(_03176_),
    .A2(_05679_),
    .B(_05681_),
    .C(_05678_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11441_ (.I(_05647_),
    .Z(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11442_ (.A1(_05480_),
    .A2(_05678_),
    .B(_05682_),
    .C(_05683_),
    .ZN(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11443_ (.I(_05659_),
    .Z(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11444_ (.I(_05663_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11445_ (.A1(_05332_),
    .A2(_05685_),
    .B1(_05686_),
    .B2(\as2650.regs[0][4] ),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11446_ (.A1(_05684_),
    .A2(_05687_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11447_ (.A1(\as2650.regs[4][5] ),
    .A2(_05680_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11448_ (.A1(_03226_),
    .A2(_05679_),
    .B(_05688_),
    .C(_05661_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11449_ (.A1(_05495_),
    .A2(_05678_),
    .B(_05689_),
    .C(_05683_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11450_ (.A1(_05336_),
    .A2(_05685_),
    .B1(_05686_),
    .B2(\as2650.regs[0][5] ),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11451_ (.A1(_05690_),
    .A2(_05691_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11452_ (.A1(\as2650.regs[4][6] ),
    .A2(_05680_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11453_ (.A1(_03268_),
    .A2(_05679_),
    .B(_05692_),
    .C(_05661_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11454_ (.A1(_05512_),
    .A2(_05678_),
    .B(_05693_),
    .C(_05683_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11455_ (.A1(_05338_),
    .A2(_05685_),
    .B1(_05686_),
    .B2(\as2650.regs[0][6] ),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11456_ (.A1(_05694_),
    .A2(_05695_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11457_ (.A1(\as2650.regs[4][7] ),
    .A2(_05680_),
    .B1(_05525_),
    .B2(_05654_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11458_ (.A1(_03315_),
    .A2(_05679_),
    .B(_05696_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11459_ (.A1(_05683_),
    .A2(_05697_),
    .ZN(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11460_ (.A1(_05340_),
    .A2(_05685_),
    .B1(_05686_),
    .B2(\as2650.regs[0][7] ),
    .ZN(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11461_ (.A1(_05698_),
    .A2(_05699_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11462_ (.A1(_02249_),
    .A2(_02420_),
    .A3(_02549_),
    .A4(_02592_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11463_ (.I(_05700_),
    .Z(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11464_ (.I0(_02548_),
    .I1(\as2650.stack[9][0] ),
    .S(_05701_),
    .Z(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11465_ (.I(_05702_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11466_ (.I0(_02553_),
    .I1(\as2650.stack[9][1] ),
    .S(_05701_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11467_ (.I(_05703_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11468_ (.I0(_02555_),
    .I1(\as2650.stack[9][2] ),
    .S(_05701_),
    .Z(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11469_ (.I(_05704_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11470_ (.I0(_02557_),
    .I1(\as2650.stack[9][3] ),
    .S(_05701_),
    .Z(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11471_ (.I(_05705_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11472_ (.I(_05700_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11473_ (.I0(_02559_),
    .I1(\as2650.stack[9][4] ),
    .S(_05706_),
    .Z(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11474_ (.I(_05707_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11475_ (.I0(_02562_),
    .I1(\as2650.stack[9][5] ),
    .S(_05706_),
    .Z(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11476_ (.I(_05708_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11477_ (.I0(_02564_),
    .I1(\as2650.stack[9][6] ),
    .S(_05706_),
    .Z(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11478_ (.I(_05709_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11479_ (.I0(_02566_),
    .I1(\as2650.stack[9][7] ),
    .S(_05706_),
    .Z(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11480_ (.I(_05710_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11481_ (.I(_05700_),
    .Z(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11482_ (.I0(_02568_),
    .I1(\as2650.stack[9][8] ),
    .S(_05711_),
    .Z(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11483_ (.I(_05712_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11484_ (.I0(_02571_),
    .I1(\as2650.stack[9][9] ),
    .S(_05711_),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11485_ (.I(_05713_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11486_ (.I0(_02573_),
    .I1(\as2650.stack[9][10] ),
    .S(_05711_),
    .Z(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11487_ (.I(_05714_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11488_ (.I0(_02575_),
    .I1(\as2650.stack[9][11] ),
    .S(_05711_),
    .Z(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11489_ (.I(_05715_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11490_ (.I(_05700_),
    .Z(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11491_ (.I0(_02577_),
    .I1(\as2650.stack[9][12] ),
    .S(_05716_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11492_ (.I(_05717_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11493_ (.I0(_02580_),
    .I1(\as2650.stack[9][13] ),
    .S(_05716_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11494_ (.I(_05718_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11495_ (.I0(_02582_),
    .I1(\as2650.stack[9][14] ),
    .S(_05716_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11496_ (.I(_05719_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11497_ (.I0(_02584_),
    .I1(\as2650.stack[9][15] ),
    .S(_05716_),
    .Z(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11498_ (.I(_05720_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11499_ (.D(_00005_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.relative_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11500_ (.D(_00006_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net114));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11501_ (.D(_00007_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net121));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11502_ (.D(_00008_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(net122));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11503_ (.D(_00009_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net123));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11504_ (.D(_00010_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(net124));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11505_ (.D(_00011_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(net125));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11506_ (.D(_00012_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(net126));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11507_ (.D(_00013_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(net127));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11508_ (.D(_00014_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(net128));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11509_ (.D(_00015_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(net129));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11510_ (.D(_00016_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(net115));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11511_ (.D(_00017_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(net116));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11512_ (.D(_00018_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(net117));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11513_ (.D(_00019_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(net118));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11514_ (.D(_00020_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(net119));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11515_ (.D(_00021_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(net120));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11516_ (.D(_00022_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(net98));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11517_ (.D(_00023_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(net105));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11518_ (.D(_00024_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(net106));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11519_ (.D(_00025_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(net107));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11520_ (.D(_00026_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(net108));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11521_ (.D(_00027_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(net109));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11522_ (.D(_00028_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(net110));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11523_ (.D(_00029_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(net111));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11524_ (.D(_00030_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(net112));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11525_ (.D(_00031_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net113));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11526_ (.D(_00032_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(net99));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11527_ (.D(_00033_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(net100));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11528_ (.D(_00034_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net101));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11529_ (.D(_00035_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(net102));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11530_ (.D(_00036_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(net103));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11531_ (.D(_00037_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(net104));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11532_ (.D(_00038_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net151));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11533_ (.D(_00039_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(net152));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11534_ (.D(_00040_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(net153));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11535_ (.D(_00041_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(net224));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11536_ (.D(_00042_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(net225));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11537_ (.D(_00043_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(net236));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11538_ (.D(_00044_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(net247));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11539_ (.D(_00045_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(net250));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11540_ (.D(_00046_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(net251));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11541_ (.D(_00047_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(net252));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11542_ (.D(_00048_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(net253));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11543_ (.D(_00049_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(net254));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11544_ (.D(_00050_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(net255));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11545_ (.D(_00051_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(net256));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11546_ (.D(_00052_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(net226));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11547_ (.D(_00053_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(net227));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11548_ (.D(_00054_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(net228));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11549_ (.D(_00055_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(net229));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11550_ (.D(_00056_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(net230));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11551_ (.D(_00057_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(net231));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11552_ (.D(_00058_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(net232));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11553_ (.D(_00059_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(net233));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11554_ (.D(_00060_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net234));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11555_ (.D(_00061_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net235));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11556_ (.D(_00062_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(net237));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11557_ (.D(_00063_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(net238));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11558_ (.D(_00064_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net239));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11559_ (.D(_00065_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(net240));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11560_ (.D(_00066_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(net241));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11561_ (.D(_00067_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(net242));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11562_ (.D(_00068_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(net243));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11563_ (.D(_00069_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(net244));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11564_ (.D(_00070_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(net245));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11565_ (.D(_00071_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(net246));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11566_ (.D(_00072_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(net248));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11567_ (.D(_00073_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(net249));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11568_ (.D(_00074_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(wb_feedback_delay));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11569_ (.D(net339),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(wb_debug_cc));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11570_ (.D(net388),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(wb_debug_carry));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11571_ (.D(net327),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\web_behavior[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11572_ (.D(net323),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\web_behavior[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11573_ (.D(net331),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(wb_reset_override_en));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11574_ (.D(net350),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(wb_reset_override));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11575_ (.D(net380),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(wb_io3_test));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11576_ (.D(net335),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(net174));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11577_ (.D(_00083_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.wb_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11578_ (.D(_00084_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\wb_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11579_ (.D(_00085_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(\wb_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11580_ (.D(_00086_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(\wb_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11581_ (.D(_00087_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\wb_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11582_ (.D(_00088_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\wb_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11583_ (.D(_00089_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\wb_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11584_ (.D(_00090_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\wb_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11585_ (.D(_00091_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\wb_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11586_ (.D(_00092_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\wb_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11587_ (.D(net366),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\wb_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11588_ (.D(net362),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\wb_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11589_ (.D(_00095_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\wb_counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11590_ (.D(net343),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\wb_counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11591_ (.D(net347),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\wb_counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11592_ (.D(net358),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\wb_counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11593_ (.D(net354),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\wb_counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11594_ (.D(_00100_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11595_ (.D(_00101_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11596_ (.D(_00102_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\wb_counter[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11597_ (.D(_00103_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\wb_counter[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11598_ (.D(_00104_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\wb_counter[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11599_ (.D(_00105_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\wb_counter[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11600_ (.D(_00106_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\wb_counter[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11601_ (.D(_00107_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\wb_counter[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11602_ (.D(_00108_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\wb_counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11603_ (.D(_00109_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\wb_counter[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11604_ (.D(_00110_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\wb_counter[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11605_ (.D(_00111_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\wb_counter[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11606_ (.D(_00112_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\wb_counter[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11607_ (.D(_00113_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\wb_counter[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11608_ (.D(_00114_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\wb_counter[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11609_ (.D(_00115_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\wb_counter[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11610_ (.D(_00116_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.chirpchar[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11611_ (.D(_00117_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11612_ (.D(_00118_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11613_ (.D(_00119_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11614_ (.D(_00120_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11615_ (.D(_00121_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11616_ (.D(_00122_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11617_ (.D(_00123_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11618_ (.D(_00124_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11619_ (.D(_00125_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11620_ (.D(_00126_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11621_ (.D(_00127_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11622_ (.D(_00128_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11623_ (.D(_00129_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11624_ (.D(_00130_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11625_ (.D(_00131_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11626_ (.D(_00132_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11627_ (.D(_00133_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11628_ (.D(_00134_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11629_ (.D(_00135_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11630_ (.D(_00136_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11631_ (.D(_00137_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11632_ (.D(_00138_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11633_ (.D(_00139_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11634_ (.D(_00140_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11635_ (.D(_00141_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11636_ (.D(_00142_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11637_ (.D(_00143_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11638_ (.D(_00144_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11639_ (.D(_00145_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00146_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11641_ (.D(_00147_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11642_ (.D(_00148_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11643_ (.D(_00149_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11644_ (.D(_00150_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11645_ (.D(_00151_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11646_ (.D(_00152_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11647_ (.D(_00153_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11648_ (.D(_00154_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11649_ (.D(_00155_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00156_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00157_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00158_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00159_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00160_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00161_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00162_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00163_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00164_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00165_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00166_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00167_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00168_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00169_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00170_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00171_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00172_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00173_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00174_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00175_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00176_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00177_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00178_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11673_ (.D(_00179_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00180_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11675_ (.D(_00000_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.chirpchar[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00001_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.chirpchar[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11677_ (.D(_00002_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.chirpchar[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00003_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.chirpchar[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11679_ (.D(_00004_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.chirpchar[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11680_ (.D(_00181_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11681_ (.D(_00182_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00183_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00184_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00185_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00186_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00187_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00188_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00189_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00190_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00191_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00192_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00193_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00194_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00195_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00196_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00197_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00198_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00199_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00200_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00201_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00202_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00203_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00204_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00205_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00206_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00207_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00208_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00209_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00210_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00211_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00212_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00213_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00214_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00215_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00216_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00217_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00218_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00219_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00220_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00221_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00222_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00223_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00224_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00225_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00226_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00227_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00228_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00229_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00230_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00231_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00232_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00233_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00234_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00235_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00236_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00237_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00238_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00239_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00240_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00241_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00242_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00243_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00244_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00245_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00246_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00247_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00248_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00249_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00250_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00251_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00252_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00253_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00254_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00255_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00256_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00257_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00258_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00259_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00260_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00261_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00262_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00263_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00264_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00265_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00266_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00267_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00268_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00269_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00270_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00271_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00272_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00273_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00274_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00275_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00276_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00277_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00278_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00279_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00280_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00281_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00282_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00283_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00284_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00285_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00286_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00287_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00288_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00289_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00290_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00291_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00292_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00293_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00294_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00295_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00296_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00297_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00298_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00299_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00300_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00301_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00302_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00303_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00304_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00305_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00306_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00307_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00308_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00309_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00310_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00311_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00312_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00313_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00314_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00315_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00316_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00317_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11817_ (.D(_00318_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00319_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00320_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00321_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00322_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00323_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00324_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00325_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00326_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00327_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00328_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00329_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00330_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00331_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00332_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00333_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00334_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00335_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00336_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00337_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00338_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00339_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00340_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11840_ (.D(_00341_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11841_ (.D(_00342_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11842_ (.D(_00343_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00344_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00345_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00346_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00347_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00348_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00349_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00350_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00351_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00352_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00353_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00354_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00355_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00356_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00357_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00358_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00359_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00360_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00361_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00362_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00363_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00364_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00365_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.last_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00366_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.last_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00367_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.last_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00368_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.last_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00369_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.last_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00370_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.last_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00371_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.last_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00372_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.last_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00373_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.chirp_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11873_ (.D(_00374_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.chirp_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00375_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.chirp_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00376_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.indirect_target[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11876_ (.D(_00377_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11877_ (.D(_00378_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00379_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.indirect_target[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00380_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.indirect_target[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00381_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.indirect_target[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00382_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.indirect_target[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00383_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.indirect_target[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00384_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.indirect_target[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00385_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.indirect_target[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00386_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.indirect_target[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00387_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.indirect_target[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00388_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00389_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00390_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00391_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.indirect_target[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11891_ (.D(_00392_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.indexed_cyc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11892_ (.D(_00393_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.indexed_cyc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00394_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.indirect_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11894_ (.D(_00395_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(net205));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11895_ (.D(_00396_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.extend ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11896_ (.D(_00397_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.warmup[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11897_ (.D(_00398_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.warmup[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00399_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00400_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00401_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00402_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.instruction_args_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00403_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.instruction_args_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00404_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.instruction_args_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00405_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.instruction_args_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00406_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.instruction_args_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11906_ (.D(_00407_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.instruction_args_latch[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00408_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.instruction_args_latch[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00409_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.instruction_args_latch[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11909_ (.D(_00410_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.instruction_args_latch[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00411_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.instruction_args_latch[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00412_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.instruction_args_latch[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11912_ (.D(_00413_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.instruction_args_latch[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00414_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.instruction_args_latch[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00415_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00416_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11916_ (.D(_00417_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11917_ (.D(_00418_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00419_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.insin[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11919_ (.D(_00420_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.insin[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00421_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.insin[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00422_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.insin[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00423_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.insin[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00424_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.insin[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11924_ (.D(_00425_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.insin[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00426_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.insin[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00427_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.page_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11927_ (.D(_00428_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.page_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00429_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.page_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11929_ (.D(_00430_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.last_addr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11930_ (.D(_00431_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.last_addr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00432_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.last_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00433_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.last_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00434_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.last_addr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00435_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.last_addr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00436_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.last_addr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00437_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.last_addr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00438_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.ivectors_base[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00439_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.ivectors_base[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00440_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.ivectors_base[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11940_ (.D(_00441_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.ivectors_base[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11941_ (.D(_00442_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.ivectors_base[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11942_ (.D(_00443_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\as2650.ivectors_base[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00444_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.ivectors_base[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_00445_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\as2650.ivectors_base[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11945_ (.D(_00446_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.ivectors_base[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00447_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.ivectors_base[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00448_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.ivectors_base[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_00449_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.ivectors_base[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_00450_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.PC[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11950_ (.D(_00451_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.PC[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11951_ (.D(_00452_),
    .CLK(clknet_4_6__leaf_wb_clk_i),
    .Q(\as2650.PC[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00453_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.PC[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00454_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.PC[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11954_ (.D(_00455_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.PC[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00456_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.PC[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11956_ (.D(_00457_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.PC[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11957_ (.D(_00458_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.PC[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00459_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.PC[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00460_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.PC[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11960_ (.D(_00461_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.PC[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11961_ (.D(_00462_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.PC[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11962_ (.D(_00463_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.debug_psl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11963_ (.D(_00464_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.debug_psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11964_ (.D(_00465_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.debug_psl[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00466_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.debug_psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00467_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.debug_psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00468_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.debug_psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00469_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_00470_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.debug_psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00471_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.debug_psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_00472_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.debug_psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_00473_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.debug_psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11973_ (.D(_00474_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.debug_psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11974_ (.D(_00475_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.debug_psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11975_ (.D(_00476_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.debug_psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11976_ (.D(_00477_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(net173));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11977_ (.D(_00478_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.debug_psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11978_ (.D(_00479_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.irqs_latch[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11979_ (.D(_00480_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.irqs_latch[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11980_ (.D(_00481_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.irqs_latch[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11981_ (.D(_00482_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.irqs_latch[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11982_ (.D(_00483_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.irqs_latch[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11983_ (.D(_00484_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.irqs_latch[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11984_ (.D(_00485_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.irqs_latch[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11985_ (.D(_00486_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.trap ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11986_ (.D(_00487_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net139));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11987_ (.D(_00488_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(net140));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11988_ (.D(_00489_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net141));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11989_ (.D(_00490_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net142));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_00491_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(net143));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_00492_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(net144));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11992_ (.D(_00493_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(net145));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_00494_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(net146));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11994_ (.D(_00495_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net138));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00496_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(net132));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_00497_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net133));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00498_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net134));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00499_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net135));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_00500_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net136));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00501_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net137));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00502_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.ext_io_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00503_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.ext_io_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12003_ (.D(_00504_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.io_bus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_00505_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.chirpchar[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12005_ (.D(_00506_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.cpu_hidden_rom_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12006_ (.D(_00507_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12007_ (.D(_00508_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12008_ (.D(_00509_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_00510_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(_00511_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_00512_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_00513_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_00514_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.regs[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(_00515_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12015_ (.D(_00516_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.regs[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12016_ (.D(_00517_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.regs[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(_00518_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.regs[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(_00519_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(_00520_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12020_ (.D(_00521_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\as2650.regs[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12021_ (.D(_00522_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.regs[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12022_ (.D(_00523_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12023_ (.D(_00524_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12024_ (.D(_00525_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12025_ (.D(_00526_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12026_ (.D(_00527_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12027_ (.D(_00528_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.regs[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12028_ (.D(_00529_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(_00530_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12030_ (.D(_00531_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12031_ (.D(_00532_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12032_ (.D(_00533_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.regs[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12033_ (.D(_00534_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12034_ (.D(_00535_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.regs[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12035_ (.D(_00536_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.regs[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(_00537_),
    .CLK(clknet_4_15__leaf_wb_clk_i),
    .Q(\as2650.regs[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_00538_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.regs[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12038_ (.D(_00539_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12039_ (.D(_00540_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.regs[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12040_ (.D(_00541_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.regs[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12041_ (.D(_00542_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\as2650.regs[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_00543_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(_00544_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(_00545_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\as2650.regs[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12045_ (.D(_00546_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(_00547_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(_00548_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12048_ (.D(_00549_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.regs[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(_00550_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.regs[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(_00551_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(_00552_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.regs[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(_00553_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12053_ (.D(_00554_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\as2650.regs[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12054_ (.D(_00555_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12055_ (.D(_00556_),
    .CLK(clknet_4_14__leaf_wb_clk_i),
    .Q(\as2650.regs[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12056_ (.D(_00557_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.regs[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12057_ (.D(_00558_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.regs[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12058_ (.D(_00559_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12059_ (.D(_00560_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12060_ (.D(_00561_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12061_ (.D(_00562_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.regs[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12062_ (.D(_00563_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12063_ (.D(_00564_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12064_ (.D(_00565_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12065_ (.D(_00566_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12066_ (.D(_00567_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12067_ (.D(_00568_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(_00569_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12069_ (.D(_00570_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12070_ (.D(_00571_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12071_ (.D(_00572_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12072_ (.D(_00573_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12073_ (.D(_00574_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12074_ (.D(_00575_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12075_ (.D(_00576_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(_00577_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12077_ (.D(_00578_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12116_ (.I(net257),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12117_ (.I(net257),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12118_ (.I(net257),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12119_ (.I(net258),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12120_ (.I(net258),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12121_ (.I(net258),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12122_ (.I(net259),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12123_ (.I(net257),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12124_ (.I(net175),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12125_ (.I(net176),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12126_ (.I(net177),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12127_ (.I(net178),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12128_ (.I(net179),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12129_ (.I(net163),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12130_ (.I(net164),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12131_ (.I(net165),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_129_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_130_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_132_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_135_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_136_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_137_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_138_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_139_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_140_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_142_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_144_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_145_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_146_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_147_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_148_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_150_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_151_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_152_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_153_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_154_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_155_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_156_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_157_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_158_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_159_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_160_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_160_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_161_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_162_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_163_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_163_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_164_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_164_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_165_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_165_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout257 (.I(net258),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout258 (.I(net156),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout259 (.I(net156),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold1 (.I(wbs_dat_i[10]),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold10 (.I(wbs_dat_i[8]),
    .Z(net421));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold100 (.I(net437),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold101 (.I(net439),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold102 (.I(net428),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold103 (.I(net438),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold104 (.I(net440),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold105 (.I(net441),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold106 (.I(net442),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold107 (.I(wbs_cyc_i),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold108 (.I(_01697_),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold109 (.I(wbs_dat_i[27]),
    .Z(net428));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold11 (.I(wbs_dat_i[4]),
    .Z(net422));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold110 (.I(wbs_dat_i[19]),
    .Z(net429));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold111 (.I(wbs_dat_i[16]),
    .Z(net430));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold112 (.I(wbs_dat_i[24]),
    .Z(net431));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold113 (.I(wbs_adr_i[19]),
    .Z(net432));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold114 (.I(wbs_dat_i[26]),
    .Z(net433));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold115 (.I(wbs_dat_i[17]),
    .Z(net434));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold116 (.I(wbs_dat_i[23]),
    .Z(net435));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold117 (.I(wbs_dat_i[22]),
    .Z(net436));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold118 (.I(wbs_dat_i[25]),
    .Z(net437));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold119 (.I(wbs_dat_i[18]),
    .Z(net438));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold12 (.I(wbs_dat_i[9]),
    .Z(net423));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold120 (.I(wbs_dat_i[31]),
    .Z(net439));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold121 (.I(wbs_dat_i[29]),
    .Z(net440));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold122 (.I(wbs_dat_i[28]),
    .Z(net441));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold123 (.I(wbs_adr_i[21]),
    .Z(net442));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold124 (.I(wbs_dat_i[11]),
    .Z(net443));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold13 (.I(wbs_dat_i[6]),
    .Z(net424));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold14 (.I(wbs_dat_i[3]),
    .Z(net425));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold15 (.I(wbs_dat_i[30]),
    .Z(net426));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold16 (.I(wbs_dat_i[21]),
    .Z(net427));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold17 (.I(net425),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold18 (.I(net89),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold19 (.I(_02000_),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold2 (.I(wbs_dat_i[20]),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold20 (.I(_00078_),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold21 (.I(net376),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold22 (.I(net86),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold23 (.I(_01998_),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold24 (.I(_00077_),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold25 (.I(net422),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold26 (.I(net90),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold27 (.I(_02003_),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold28 (.I(_00079_),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold29 (.I(net419),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold3 (.I(wbs_dat_i[1]),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold30 (.I(net93),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold31 (.I(_02008_),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold32 (.I(_00082_),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold33 (.I(net420),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold34 (.I(net64),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold35 (.I(_01991_),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold36 (.I(_00075_),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold37 (.I(net390),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold38 (.I(net67),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold39 (.I(_02066_),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold4 (.I(wbs_dat_i[5]),
    .Z(net415));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold40 (.I(_00096_),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold41 (.I(net389),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold42 (.I(net68),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold43 (.I(_02068_),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold44 (.I(_00097_),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold45 (.I(net415),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold46 (.I(_02005_),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold47 (.I(_00080_),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold48 (.I(wbs_dat_i[15]),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold49 (.I(net70),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold5 (.I(wbs_adr_i[22]),
    .Z(net416));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold50 (.I(_02079_),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold51 (.I(_00099_),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold52 (.I(net392),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold53 (.I(net69),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold54 (.I(_02071_),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold55 (.I(_00098_),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold56 (.I(net412),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold57 (.I(net65),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold58 (.I(_02055_),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold59 (.I(_00094_),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold6 (.I(_01919_),
    .Z(net417));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold60 (.I(net423),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold61 (.I(net95),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold62 (.I(_02052_),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold63 (.I(_00093_),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold64 (.I(net416),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold65 (.I(_02012_),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold66 (.I(net443),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold67 (.I(net66),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold68 (.I(net421),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold69 (.I(net94),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold7 (.I(_01987_),
    .Z(net418));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold70 (.I(net430),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold71 (.I(net71),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold72 (.I(_01727_),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold73 (.I(wbs_dat_i[2]),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold74 (.I(net424),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold75 (.I(net92),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold76 (.I(_02007_),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold77 (.I(_00081_),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold78 (.I(wbs_adr_i[20]),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold79 (.I(_01701_),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold8 (.I(wbs_dat_i[7]),
    .Z(net419));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold80 (.I(_01702_),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold81 (.I(_01703_),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold82 (.I(_01724_),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold83 (.I(net414),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold84 (.I(_01995_),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold85 (.I(_00076_),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold86 (.I(wbs_dat_i[13]),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold87 (.I(wbs_dat_i[12]),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold88 (.I(net413),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold89 (.I(wbs_dat_i[14]),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold9 (.I(wbs_dat_i[0]),
    .Z(net420));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold90 (.I(net429),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold91 (.I(net427),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold92 (.I(net431),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold93 (.I(net436),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold94 (.I(net433),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold95 (.I(net435),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold96 (.I(net426),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold97 (.I(net432),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 hold98 (.I(_01753_),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 hold99 (.I(net434),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(bus_in_gpios[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(bus_in_serial_ports[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(bus_in_serial_ports[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(bus_in_serial_ports[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(bus_in_serial_ports[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(bus_in_serial_ports[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(bus_in_serial_ports[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(bus_in_serial_ports[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(bus_in_sid[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(bus_in_sid[1]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(bus_in_sid[2]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(bus_in_gpios[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(bus_in_sid[3]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(bus_in_sid[4]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(bus_in_sid[5]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(bus_in_sid[6]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(bus_in_sid[7]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(bus_in_timers[0]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(bus_in_timers[1]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(bus_in_timers[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(bus_in_timers[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(bus_in_timers[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(bus_in_gpios[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(bus_in_timers[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(bus_in_timers[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(bus_in_timers[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input33 (.I(io_in[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input34 (.I(io_in[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input35 (.I(io_in[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input36 (.I(io_in[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input37 (.I(io_in[4]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input38 (.I(io_in[5]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input39 (.I(io_in[6]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(bus_in_gpios[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input40 (.I(io_in[7]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input41 (.I(io_in[8]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input42 (.I(io_in[9]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input43 (.I(irqs[0]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input44 (.I(irqs[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input45 (.I(irqs[2]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(irqs[3]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input47 (.I(irqs[4]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input48 (.I(irqs[5]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(irqs[6]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(bus_in_gpios[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input50 (.I(rom_bus_in[0]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input51 (.I(rom_bus_in[1]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input52 (.I(rom_bus_in[2]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input53 (.I(rom_bus_in[3]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input54 (.I(rom_bus_in[4]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input55 (.I(rom_bus_in[5]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input56 (.I(rom_bus_in[6]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input57 (.I(rom_bus_in[7]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input58 (.I(wb_rst_i),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input59 (.I(net400),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(bus_in_gpios[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input60 (.I(net381),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input61 (.I(net409),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input62 (.I(net367),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(net410),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input64 (.I(net336),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(net359),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(net369),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(net340),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(net344),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(net355),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(bus_in_gpios[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(net351),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(net373),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(net402),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(net406),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(net393),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input75 (.I(net386),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(net391),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(net394),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(net396),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(net398),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(bus_in_gpios[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(net395),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input81 (.I(net403),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input82 (.I(net397),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input83 (.I(net405),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input84 (.I(net408),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input85 (.I(net407),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input86 (.I(net324),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input87 (.I(net399),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input88 (.I(net404),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(net320),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(bus_in_serial_ports[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input90 (.I(net328),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input91 (.I(net348),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input92 (.I(net377),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input93 (.I(net332),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input94 (.I(net371),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input95 (.I(net363),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input96 (.I(wbs_stb_i),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input97 (.I(wbs_we_i),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap260 (.I(_01432_),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap262 (.I(net263),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 max_cap264 (.I(_00942_),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output100 (.I(net100),
    .Z(RAM_end_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output101 (.I(net101),
    .Z(RAM_end_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output102 (.I(net102),
    .Z(RAM_end_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output103 (.I(net103),
    .Z(RAM_end_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output104 (.I(net104),
    .Z(RAM_end_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output105 (.I(net105),
    .Z(RAM_end_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(RAM_end_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(RAM_end_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(RAM_end_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(RAM_end_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(RAM_end_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(RAM_end_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(RAM_end_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(RAM_end_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(RAM_start_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(RAM_start_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(RAM_start_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(RAM_start_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(RAM_start_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(RAM_start_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(RAM_start_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(RAM_start_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(RAM_start_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(RAM_start_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(RAM_start_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(RAM_start_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output126 (.I(net126),
    .Z(RAM_start_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output127 (.I(net127),
    .Z(RAM_start_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output128 (.I(net128),
    .Z(RAM_start_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output129 (.I(net129),
    .Z(RAM_start_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output130 (.I(net130),
    .Z(WEb_raw));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output131 (.I(net131),
    .Z(boot_rom_en));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output132 (.I(net132),
    .Z(bus_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output133 (.I(net133),
    .Z(bus_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output134 (.I(net134),
    .Z(bus_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output135 (.I(net135),
    .Z(bus_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output136 (.I(net136),
    .Z(bus_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output137 (.I(net137),
    .Z(bus_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output138 (.I(net138),
    .Z(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output139 (.I(net139),
    .Z(bus_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output140 (.I(net140),
    .Z(bus_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output141 (.I(net141),
    .Z(bus_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output142 (.I(net142),
    .Z(bus_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output143 (.I(net143),
    .Z(bus_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output144 (.I(net144),
    .Z(bus_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output145 (.I(net145),
    .Z(bus_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output146 (.I(net146),
    .Z(bus_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output147 (.I(net147),
    .Z(bus_we_gpios));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output148 (.I(net148),
    .Z(bus_we_serial_ports));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output149 (.I(net149),
    .Z(bus_we_sid));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output150 (.I(net150),
    .Z(bus_we_timers));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output151 (.I(net151),
    .Z(cs_port[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output152 (.I(net152),
    .Z(cs_port[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output153 (.I(net153),
    .Z(cs_port[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output154 (.I(net154),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output155 (.I(net155),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output156 (.I(net259),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output157 (.I(net157),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output158 (.I(net158),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output159 (.I(net159),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output160 (.I(net160),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output161 (.I(net161),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output162 (.I(net162),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output163 (.I(net163),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output164 (.I(net164),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output165 (.I(net165),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output166 (.I(net166),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output167 (.I(net167),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output168 (.I(net168),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output169 (.I(net169),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output170 (.I(net170),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output171 (.I(net171),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output172 (.I(net172),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output173 (.I(net173),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output174 (.I(net174),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output175 (.I(net175),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output176 (.I(net176),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output177 (.I(net177),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output178 (.I(net178),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output179 (.I(net179),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output180 (.I(net180),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output181 (.I(net181),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output182 (.I(net182),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output183 (.I(net183),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output184 (.I(net184),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output185 (.I(net185),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output186 (.I(net186),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output187 (.I(net187),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output188 (.I(net188),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output189 (.I(net189),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output190 (.I(net190),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output191 (.I(net191),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output192 (.I(net192),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output193 (.I(net193),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output194 (.I(net194),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output195 (.I(net195),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output196 (.I(net196),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output197 (.I(net197),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output198 (.I(net198),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output199 (.I(net199),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output200 (.I(net200),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output201 (.I(net201),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output202 (.I(net202),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output203 (.I(net203),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output204 (.I(net204),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output205 (.I(net205),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output206 (.I(net206),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output207 (.I(net207),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output208 (.I(net208),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output209 (.I(net209),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output210 (.I(net210),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output211 (.I(net211),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output212 (.I(net212),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output213 (.I(net213),
    .Z(le_hi_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output214 (.I(net214),
    .Z(le_lo_act));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output215 (.I(net215),
    .Z(reset_out));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output216 (.I(net216),
    .Z(rom_bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output217 (.I(net217),
    .Z(rom_bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output218 (.I(net218),
    .Z(rom_bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output219 (.I(net219),
    .Z(rom_bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output220 (.I(net220),
    .Z(rom_bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output221 (.I(net221),
    .Z(rom_bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output222 (.I(net222),
    .Z(rom_bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output223 (.I(net223),
    .Z(rom_bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output224 (.I(net224),
    .Z(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output225 (.I(net225),
    .Z(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output226 (.I(net226),
    .Z(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output227 (.I(net227),
    .Z(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output228 (.I(net228),
    .Z(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output229 (.I(net229),
    .Z(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output230 (.I(net230),
    .Z(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output231 (.I(net231),
    .Z(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output232 (.I(net232),
    .Z(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output233 (.I(net233),
    .Z(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output234 (.I(net234),
    .Z(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output235 (.I(net235),
    .Z(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output236 (.I(net236),
    .Z(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output237 (.I(net237),
    .Z(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output238 (.I(net238),
    .Z(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output239 (.I(net239),
    .Z(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output240 (.I(net240),
    .Z(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output241 (.I(net241),
    .Z(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output242 (.I(net242),
    .Z(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output243 (.I(net243),
    .Z(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output244 (.I(net244),
    .Z(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output245 (.I(net245),
    .Z(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output246 (.I(net246),
    .Z(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output247 (.I(net247),
    .Z(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output248 (.I(net248),
    .Z(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output249 (.I(net249),
    .Z(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output250 (.I(net250),
    .Z(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output251 (.I(net251),
    .Z(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output252 (.I(net252),
    .Z(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output253 (.I(net253),
    .Z(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output254 (.I(net254),
    .Z(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output255 (.I(net255),
    .Z(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output256 (.I(net256),
    .Z(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output98 (.I(net98),
    .Z(RAM_end_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output99 (.I(net99),
    .Z(RAM_end_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 rebuffer1 (.I(_00776_),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer10 (.I(_00767_),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer11 (.I(_01110_),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer12 (.I(_03491_),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 rebuffer13 (.I(_00776_),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer14 (.I(_00889_),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer15 (.I(\as2650.cycle[3] ),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer16 (.I(\as2650.cycle[2] ),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer2 (.I(net304),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer3 (.I(net304),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 rebuffer4 (.I(_00785_),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_01112_),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer6 (.I(_01031_),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer7 (.I(_00767_),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer8 (.I(_00891_),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 rebuffer9 (.I(net311),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire261 (.I(net263),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire263 (.I(_04799_),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_286 (.Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_287 (.Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_288 (.Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_289 (.Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_290 (.Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_291 (.Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_292 (.Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_293 (.Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_294 (.Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_295 (.Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_296 (.Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_297 (.Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_298 (.Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_299 (.Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_300 (.Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_301 (.Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_302 (.Z(net302));
 assign io_oeb[0] = net286;
 assign io_oeb[13] = net267;
 assign io_oeb[14] = net268;
 assign io_oeb[15] = net269;
 assign io_oeb[16] = net270;
 assign io_oeb[17] = net271;
 assign io_oeb[18] = net272;
 assign io_oeb[1] = net265;
 assign io_oeb[2] = net266;
 assign io_oeb[4] = net287;
 assign io_out[0] = net273;
 assign io_out[4] = net274;
 assign irq[0] = net275;
 assign irq[1] = net276;
 assign irq[2] = net277;
 assign la_data_out[33] = net288;
 assign la_data_out[34] = net289;
 assign la_data_out[35] = net290;
 assign la_data_out[36] = net291;
 assign la_data_out[37] = net292;
 assign la_data_out[38] = net293;
 assign la_data_out[39] = net294;
 assign la_data_out[40] = net295;
 assign la_data_out[41] = net278;
 assign la_data_out[42] = net279;
 assign la_data_out[43] = net280;
 assign la_data_out[44] = net281;
 assign la_data_out[45] = net282;
 assign la_data_out[46] = net283;
 assign la_data_out[47] = net284;
 assign la_data_out[48] = net285;
 assign la_data_out[49] = net296;
 assign la_data_out[50] = net297;
 assign la_data_out[51] = net298;
 assign la_data_out[52] = net299;
 assign la_data_out[53] = net300;
 assign la_data_out[54] = net301;
 assign la_data_out[55] = net302;
endmodule

